* NGSPICE file created from bias_cell.ext - technology: sky130A

X0 BIAS1 ADC_ON BIAS1_OUT GND sky130_fd_pr__nfet_01v8 ad=2.5e+12p pd=1.1e+07u as=5.9425e+12p ps=1.514e+07u w=5e+06u l=1e+06u
X1 NB1 NB1 GND GND sky130_fd_pr__nfet_01v8_lvt ad=3.5e+11p pd=2.7e+06u as=1.237e+13p ps=4.654e+07u w=1e+06u l=1.2e+06u
X2 BIAS2_OUT BIAS2_OUT GND GND sky130_fd_pr__nfet_01v8_lvt ad=5.9725e+12p pd=1.52e+07u as=0p ps=0u w=1e+06u l=1e+06u
X3 NB2 NB2 GND GND sky130_fd_pr__nfet_01v8_lvt ad=3.5e+11p pd=2.7e+06u as=0p ps=0u w=1e+06u l=1.2e+06u
X4 BIAS2 ADC_ON BIAS2_OUT GND sky130_fd_pr__nfet_01v8 ad=2.5e+12p pd=1.1e+07u as=0p ps=0u w=5e+06u l=1e+06u
X5 AMP_IB AMP_IB GND GND sky130_fd_pr__nfet_01v8_lvt ad=5.6e+12p pd=1.74e+07u as=0p ps=0u w=8e+06u l=2e+06u
X6 OUT_IB OUT_IB GND GND sky130_fd_pr__nfet_01v8_lvt ad=5.6e+12p pd=1.74e+07u as=0p ps=0u w=8e+06u l=2e+06u
X7 BIAS1_OUT BIAS1_OUT GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X8 SF_IB SF_IB VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=5.5e+11p pd=3.1e+06u as=4.5e+11p ps=2.9e+06u w=1e+06u l=1e+06u
.end
