magic
tech sky130B
magscale 1 2
timestamp 1608136834
<< nwell >>
rect 56024 -71632 85570 -69172
rect 64460 -72444 65422 -72442
rect 56156 -88598 65422 -72444
rect 78152 -72919 85563 -71632
rect 78152 -72934 84340 -72919
rect 56156 -88602 64500 -88598
<< pwell >>
rect 65600 -88466 86317 -87472
rect 65600 -89064 86349 -88466
rect 54937 -89070 86349 -89064
rect 54937 -89072 68152 -89070
rect 54937 -89074 66544 -89072
rect 66866 -89074 66900 -89072
rect 67222 -89074 67256 -89072
rect 68330 -89074 86349 -89070
rect 54937 -90229 86349 -89074
rect 54937 -91879 86351 -90229
<< psubdiff >>
rect 54994 -91166 86026 -91122
rect 54994 -91200 55128 -91166
rect 85920 -91200 86026 -91166
rect 54994 -91240 86026 -91200
rect 54994 -91274 55130 -91240
rect 85922 -91274 86026 -91240
rect 54994 -91314 86026 -91274
rect 54994 -91348 55132 -91314
rect 85924 -91348 86026 -91314
rect 54994 -91388 86026 -91348
rect 54994 -91422 55134 -91388
rect 85926 -91422 86026 -91388
rect 54994 -91462 86026 -91422
rect 54994 -91496 55136 -91462
rect 85928 -91496 86026 -91462
rect 54994 -91536 86026 -91496
rect 54994 -91570 55136 -91536
rect 85928 -91570 86026 -91536
rect 54994 -91610 86026 -91570
rect 54994 -91644 55138 -91610
rect 85930 -91644 86026 -91610
rect 54994 -91684 86026 -91644
rect 54994 -91718 55136 -91684
rect 85928 -91718 86026 -91684
rect 54994 -91758 86026 -91718
rect 54994 -91792 55148 -91758
rect 85940 -91792 86026 -91758
rect 54994 -91832 86026 -91792
rect 54994 -91866 55146 -91832
rect 85938 -91866 86026 -91832
rect 54994 -91898 86026 -91866
<< nsubdiff >>
rect 56126 -69352 83544 -69350
rect 56126 -69396 84298 -69352
rect 56126 -69430 69062 -69396
rect 83378 -69430 84298 -69396
rect 56126 -69434 84298 -69430
rect 56126 -69468 56212 -69434
rect 64732 -69468 84298 -69434
rect 56126 -69470 84298 -69468
rect 56126 -69504 69064 -69470
rect 83380 -69504 84298 -69470
rect 56126 -69508 84298 -69504
rect 56126 -69542 56208 -69508
rect 64728 -69542 84298 -69508
rect 56126 -69544 84298 -69542
rect 56126 -69578 69068 -69544
rect 83384 -69578 84298 -69544
rect 56126 -69582 84298 -69578
rect 56126 -69616 56208 -69582
rect 64728 -69616 84298 -69582
rect 56126 -69618 84298 -69616
rect 56126 -69652 69072 -69618
rect 83388 -69652 84298 -69618
rect 56126 -69656 84298 -69652
rect 56126 -69690 56206 -69656
rect 64726 -69690 84298 -69656
rect 56126 -69924 84298 -69690
rect 56152 -69926 84298 -69924
rect 56192 -69934 84298 -69926
rect 56260 -76560 56294 -76524
rect 64214 -76560 64282 -76524
rect 56258 -76712 56296 -76674
rect 64212 -76712 64286 -76674
rect 56268 -80546 56300 -80506
rect 64204 -80546 64298 -80506
rect 56264 -80698 56296 -80658
rect 64218 -80698 64294 -80658
rect 56238 -84402 56294 -84362
rect 64212 -84402 64268 -84362
rect 56246 -84546 56294 -84508
rect 64196 -84546 64276 -84508
rect 56334 -88100 56390 -88060
rect 64308 -88100 64364 -88060
rect 56342 -88244 56390 -88206
rect 64292 -88244 64372 -88206
<< psubdiffcont >>
rect 55128 -91200 85920 -91166
rect 55130 -91274 85922 -91240
rect 55132 -91348 85924 -91314
rect 55134 -91422 85926 -91388
rect 55136 -91496 85928 -91462
rect 55136 -91570 85928 -91536
rect 55138 -91644 85930 -91610
rect 55136 -91718 85928 -91684
rect 55148 -91792 85940 -91758
rect 55146 -91866 85938 -91832
<< nsubdiffcont >>
rect 69062 -69430 83378 -69396
rect 56212 -69468 64732 -69434
rect 69064 -69504 83380 -69470
rect 56208 -69542 64728 -69508
rect 69068 -69578 83384 -69544
rect 56208 -69616 64728 -69582
rect 69072 -69652 83388 -69618
rect 56206 -69690 64726 -69656
rect 56294 -76560 64214 -76524
rect 56296 -76712 64212 -76674
rect 56300 -80546 64204 -80506
rect 56296 -80698 64218 -80658
rect 56294 -84402 64212 -84362
rect 56294 -84546 64196 -84508
rect 56390 -88100 64308 -88060
rect 56390 -88244 64292 -88206
<< locali >>
rect 56260 -76560 56294 -76524
rect 64214 -76560 64282 -76524
rect 56258 -76712 56296 -76674
rect 64212 -76712 64286 -76674
rect 56268 -80546 56300 -80506
rect 64204 -80546 64298 -80506
rect 56264 -80698 56296 -80658
rect 64218 -80698 64294 -80658
rect 56238 -84402 56294 -84362
rect 64212 -84402 64268 -84362
rect 56246 -84546 56294 -84508
rect 64196 -84546 64276 -84508
rect 56334 -88100 56390 -88060
rect 64308 -88100 64364 -88060
rect 56392 -88168 56400 -88134
rect 56434 -88168 56472 -88134
rect 56506 -88168 56544 -88134
rect 56578 -88168 56616 -88134
rect 56650 -88168 56688 -88134
rect 56722 -88168 56760 -88134
rect 56794 -88168 56832 -88134
rect 56866 -88168 56904 -88134
rect 56938 -88168 56976 -88134
rect 57010 -88168 57048 -88134
rect 57082 -88168 57120 -88134
rect 57154 -88168 57192 -88134
rect 57226 -88168 57264 -88134
rect 57298 -88168 57336 -88134
rect 57370 -88168 57408 -88134
rect 57442 -88168 57480 -88134
rect 57514 -88168 57552 -88134
rect 57586 -88168 57624 -88134
rect 57658 -88168 57696 -88134
rect 57730 -88168 57768 -88134
rect 57802 -88168 57840 -88134
rect 57874 -88168 57912 -88134
rect 57946 -88168 57984 -88134
rect 58018 -88168 58056 -88134
rect 58090 -88168 58128 -88134
rect 58162 -88168 58200 -88134
rect 58234 -88168 58272 -88134
rect 58306 -88168 58344 -88134
rect 58378 -88168 58416 -88134
rect 58450 -88168 58488 -88134
rect 58522 -88168 58560 -88134
rect 58594 -88168 58632 -88134
rect 58666 -88168 58704 -88134
rect 58738 -88168 58776 -88134
rect 58810 -88168 58848 -88134
rect 58882 -88168 58920 -88134
rect 58954 -88168 58992 -88134
rect 59026 -88168 59064 -88134
rect 59098 -88168 59136 -88134
rect 59170 -88168 59208 -88134
rect 59242 -88168 59280 -88134
rect 59314 -88168 59352 -88134
rect 59386 -88168 59424 -88134
rect 59458 -88168 59496 -88134
rect 59530 -88168 59568 -88134
rect 59602 -88168 59640 -88134
rect 59674 -88168 59712 -88134
rect 59746 -88168 59784 -88134
rect 59818 -88168 59856 -88134
rect 59890 -88168 59928 -88134
rect 59962 -88168 60000 -88134
rect 60034 -88168 60072 -88134
rect 60106 -88168 60144 -88134
rect 60178 -88168 60216 -88134
rect 60250 -88168 60288 -88134
rect 60322 -88168 60360 -88134
rect 60394 -88168 60432 -88134
rect 60466 -88168 60504 -88134
rect 60538 -88168 60576 -88134
rect 60610 -88168 60648 -88134
rect 60682 -88168 60720 -88134
rect 60754 -88168 60792 -88134
rect 60826 -88168 60864 -88134
rect 60898 -88168 60936 -88134
rect 60970 -88168 61008 -88134
rect 61042 -88168 61080 -88134
rect 61114 -88168 61152 -88134
rect 61186 -88168 61224 -88134
rect 61258 -88168 61296 -88134
rect 61330 -88168 61368 -88134
rect 61402 -88168 61440 -88134
rect 61474 -88168 61512 -88134
rect 61546 -88168 61584 -88134
rect 61618 -88168 61656 -88134
rect 61690 -88168 61728 -88134
rect 61762 -88168 61800 -88134
rect 61834 -88168 61872 -88134
rect 61906 -88168 61944 -88134
rect 61978 -88168 62016 -88134
rect 62050 -88168 62088 -88134
rect 62122 -88168 62160 -88134
rect 62194 -88168 62232 -88134
rect 62266 -88168 62304 -88134
rect 62338 -88168 62376 -88134
rect 62410 -88168 62448 -88134
rect 62482 -88168 62520 -88134
rect 62554 -88168 62592 -88134
rect 62626 -88168 62664 -88134
rect 62698 -88168 62736 -88134
rect 62770 -88168 62808 -88134
rect 62842 -88168 62880 -88134
rect 62914 -88168 62952 -88134
rect 62986 -88168 63024 -88134
rect 63058 -88168 63096 -88134
rect 63130 -88168 63168 -88134
rect 63202 -88168 63240 -88134
rect 63274 -88168 63312 -88134
rect 63346 -88168 63384 -88134
rect 63418 -88168 63456 -88134
rect 63490 -88168 63528 -88134
rect 63562 -88168 63600 -88134
rect 63634 -88168 63672 -88134
rect 63706 -88168 63744 -88134
rect 63778 -88168 63816 -88134
rect 63850 -88168 63888 -88134
rect 63922 -88168 63960 -88134
rect 63994 -88168 64032 -88134
rect 64066 -88168 64104 -88134
rect 64138 -88168 64176 -88134
rect 64210 -88168 64248 -88134
rect 64282 -88168 64312 -88134
rect 56342 -88244 56390 -88206
rect 64292 -88244 64372 -88206
<< viali >>
rect 56400 -88094 56434 -88060
rect 56472 -88094 56506 -88060
rect 56544 -88094 56578 -88060
rect 56616 -88094 56650 -88060
rect 56688 -88094 56722 -88060
rect 56760 -88094 56794 -88060
rect 56832 -88094 56866 -88060
rect 56904 -88094 56938 -88060
rect 56976 -88094 57010 -88060
rect 57048 -88094 57082 -88060
rect 57120 -88094 57154 -88060
rect 57192 -88094 57226 -88060
rect 57264 -88094 57298 -88060
rect 57336 -88094 57370 -88060
rect 57408 -88094 57442 -88060
rect 57480 -88094 57514 -88060
rect 57552 -88094 57586 -88060
rect 57624 -88094 57658 -88060
rect 57696 -88094 57730 -88060
rect 57768 -88094 57802 -88060
rect 57840 -88094 57874 -88060
rect 57912 -88094 57946 -88060
rect 57984 -88094 58018 -88060
rect 58056 -88094 58090 -88060
rect 58128 -88094 58162 -88060
rect 58200 -88094 58234 -88060
rect 58272 -88094 58306 -88060
rect 58344 -88094 58378 -88060
rect 58416 -88094 58450 -88060
rect 58488 -88094 58522 -88060
rect 58560 -88094 58594 -88060
rect 58632 -88094 58666 -88060
rect 58704 -88094 58738 -88060
rect 58776 -88094 58810 -88060
rect 58848 -88094 58882 -88060
rect 58920 -88094 58954 -88060
rect 58992 -88094 59026 -88060
rect 59064 -88094 59098 -88060
rect 59136 -88094 59170 -88060
rect 59208 -88094 59242 -88060
rect 59280 -88094 59314 -88060
rect 59352 -88094 59386 -88060
rect 59424 -88094 59458 -88060
rect 59496 -88094 59530 -88060
rect 59568 -88094 59602 -88060
rect 59640 -88094 59674 -88060
rect 59712 -88094 59746 -88060
rect 59784 -88094 59818 -88060
rect 59856 -88094 59890 -88060
rect 59928 -88094 59962 -88060
rect 60000 -88094 60034 -88060
rect 60072 -88094 60106 -88060
rect 60144 -88094 60178 -88060
rect 60216 -88094 60250 -88060
rect 60288 -88094 60322 -88060
rect 60360 -88094 60394 -88060
rect 60432 -88094 60466 -88060
rect 60504 -88094 60538 -88060
rect 60576 -88094 60610 -88060
rect 60648 -88094 60682 -88060
rect 60720 -88094 60754 -88060
rect 60792 -88094 60826 -88060
rect 60864 -88094 60898 -88060
rect 60936 -88094 60970 -88060
rect 61008 -88094 61042 -88060
rect 61080 -88094 61114 -88060
rect 61152 -88094 61186 -88060
rect 61224 -88094 61258 -88060
rect 61296 -88094 61330 -88060
rect 61368 -88094 61402 -88060
rect 61440 -88094 61474 -88060
rect 61512 -88094 61546 -88060
rect 61584 -88094 61618 -88060
rect 61656 -88094 61690 -88060
rect 61728 -88094 61762 -88060
rect 61800 -88094 61834 -88060
rect 61872 -88094 61906 -88060
rect 61944 -88094 61978 -88060
rect 62016 -88094 62050 -88060
rect 62088 -88094 62122 -88060
rect 62160 -88094 62194 -88060
rect 62232 -88094 62266 -88060
rect 62304 -88094 62338 -88060
rect 62376 -88094 62410 -88060
rect 62448 -88094 62482 -88060
rect 62520 -88094 62554 -88060
rect 62592 -88094 62626 -88060
rect 62664 -88094 62698 -88060
rect 62736 -88094 62770 -88060
rect 62808 -88094 62842 -88060
rect 62880 -88094 62914 -88060
rect 62952 -88094 62986 -88060
rect 63024 -88094 63058 -88060
rect 63096 -88094 63130 -88060
rect 63168 -88094 63202 -88060
rect 63240 -88094 63274 -88060
rect 63312 -88094 63346 -88060
rect 63384 -88094 63418 -88060
rect 63456 -88094 63490 -88060
rect 63528 -88094 63562 -88060
rect 63600 -88094 63634 -88060
rect 63672 -88094 63706 -88060
rect 63744 -88094 63778 -88060
rect 63816 -88094 63850 -88060
rect 63888 -88094 63922 -88060
rect 63960 -88094 63994 -88060
rect 64032 -88094 64066 -88060
rect 64104 -88094 64138 -88060
rect 64176 -88094 64210 -88060
rect 64248 -88094 64282 -88060
rect 56400 -88168 56434 -88134
rect 56472 -88168 56506 -88134
rect 56544 -88168 56578 -88134
rect 56616 -88168 56650 -88134
rect 56688 -88168 56722 -88134
rect 56760 -88168 56794 -88134
rect 56832 -88168 56866 -88134
rect 56904 -88168 56938 -88134
rect 56976 -88168 57010 -88134
rect 57048 -88168 57082 -88134
rect 57120 -88168 57154 -88134
rect 57192 -88168 57226 -88134
rect 57264 -88168 57298 -88134
rect 57336 -88168 57370 -88134
rect 57408 -88168 57442 -88134
rect 57480 -88168 57514 -88134
rect 57552 -88168 57586 -88134
rect 57624 -88168 57658 -88134
rect 57696 -88168 57730 -88134
rect 57768 -88168 57802 -88134
rect 57840 -88168 57874 -88134
rect 57912 -88168 57946 -88134
rect 57984 -88168 58018 -88134
rect 58056 -88168 58090 -88134
rect 58128 -88168 58162 -88134
rect 58200 -88168 58234 -88134
rect 58272 -88168 58306 -88134
rect 58344 -88168 58378 -88134
rect 58416 -88168 58450 -88134
rect 58488 -88168 58522 -88134
rect 58560 -88168 58594 -88134
rect 58632 -88168 58666 -88134
rect 58704 -88168 58738 -88134
rect 58776 -88168 58810 -88134
rect 58848 -88168 58882 -88134
rect 58920 -88168 58954 -88134
rect 58992 -88168 59026 -88134
rect 59064 -88168 59098 -88134
rect 59136 -88168 59170 -88134
rect 59208 -88168 59242 -88134
rect 59280 -88168 59314 -88134
rect 59352 -88168 59386 -88134
rect 59424 -88168 59458 -88134
rect 59496 -88168 59530 -88134
rect 59568 -88168 59602 -88134
rect 59640 -88168 59674 -88134
rect 59712 -88168 59746 -88134
rect 59784 -88168 59818 -88134
rect 59856 -88168 59890 -88134
rect 59928 -88168 59962 -88134
rect 60000 -88168 60034 -88134
rect 60072 -88168 60106 -88134
rect 60144 -88168 60178 -88134
rect 60216 -88168 60250 -88134
rect 60288 -88168 60322 -88134
rect 60360 -88168 60394 -88134
rect 60432 -88168 60466 -88134
rect 60504 -88168 60538 -88134
rect 60576 -88168 60610 -88134
rect 60648 -88168 60682 -88134
rect 60720 -88168 60754 -88134
rect 60792 -88168 60826 -88134
rect 60864 -88168 60898 -88134
rect 60936 -88168 60970 -88134
rect 61008 -88168 61042 -88134
rect 61080 -88168 61114 -88134
rect 61152 -88168 61186 -88134
rect 61224 -88168 61258 -88134
rect 61296 -88168 61330 -88134
rect 61368 -88168 61402 -88134
rect 61440 -88168 61474 -88134
rect 61512 -88168 61546 -88134
rect 61584 -88168 61618 -88134
rect 61656 -88168 61690 -88134
rect 61728 -88168 61762 -88134
rect 61800 -88168 61834 -88134
rect 61872 -88168 61906 -88134
rect 61944 -88168 61978 -88134
rect 62016 -88168 62050 -88134
rect 62088 -88168 62122 -88134
rect 62160 -88168 62194 -88134
rect 62232 -88168 62266 -88134
rect 62304 -88168 62338 -88134
rect 62376 -88168 62410 -88134
rect 62448 -88168 62482 -88134
rect 62520 -88168 62554 -88134
rect 62592 -88168 62626 -88134
rect 62664 -88168 62698 -88134
rect 62736 -88168 62770 -88134
rect 62808 -88168 62842 -88134
rect 62880 -88168 62914 -88134
rect 62952 -88168 62986 -88134
rect 63024 -88168 63058 -88134
rect 63096 -88168 63130 -88134
rect 63168 -88168 63202 -88134
rect 63240 -88168 63274 -88134
rect 63312 -88168 63346 -88134
rect 63384 -88168 63418 -88134
rect 63456 -88168 63490 -88134
rect 63528 -88168 63562 -88134
rect 63600 -88168 63634 -88134
rect 63672 -88168 63706 -88134
rect 63744 -88168 63778 -88134
rect 63816 -88168 63850 -88134
rect 63888 -88168 63922 -88134
rect 63960 -88168 63994 -88134
rect 64032 -88168 64066 -88134
rect 64104 -88168 64138 -88134
rect 64176 -88168 64210 -88134
rect 64248 -88168 64282 -88134
rect 56400 -88242 56434 -88208
rect 56472 -88242 56506 -88208
rect 56544 -88242 56578 -88208
rect 56616 -88242 56650 -88208
rect 56688 -88242 56722 -88208
rect 56760 -88242 56794 -88208
rect 56832 -88242 56866 -88208
rect 56904 -88242 56938 -88208
rect 56976 -88242 57010 -88208
rect 57048 -88242 57082 -88208
rect 57120 -88242 57154 -88208
rect 57192 -88242 57226 -88208
rect 57264 -88242 57298 -88208
rect 57336 -88242 57370 -88208
rect 57408 -88242 57442 -88208
rect 57480 -88242 57514 -88208
rect 57552 -88242 57586 -88208
rect 57624 -88242 57658 -88208
rect 57696 -88242 57730 -88208
rect 57768 -88242 57802 -88208
rect 57840 -88242 57874 -88208
rect 57912 -88242 57946 -88208
rect 57984 -88242 58018 -88208
rect 58056 -88242 58090 -88208
rect 58128 -88242 58162 -88208
rect 58200 -88242 58234 -88208
rect 58272 -88242 58306 -88208
rect 58344 -88242 58378 -88208
rect 58416 -88242 58450 -88208
rect 58488 -88242 58522 -88208
rect 58560 -88242 58594 -88208
rect 58632 -88242 58666 -88208
rect 58704 -88242 58738 -88208
rect 58776 -88242 58810 -88208
rect 58848 -88242 58882 -88208
rect 58920 -88242 58954 -88208
rect 58992 -88242 59026 -88208
rect 59064 -88242 59098 -88208
rect 59136 -88242 59170 -88208
rect 59208 -88242 59242 -88208
rect 59280 -88242 59314 -88208
rect 59352 -88242 59386 -88208
rect 59424 -88242 59458 -88208
rect 59496 -88242 59530 -88208
rect 59568 -88242 59602 -88208
rect 59640 -88242 59674 -88208
rect 59712 -88242 59746 -88208
rect 59784 -88242 59818 -88208
rect 59856 -88242 59890 -88208
rect 59928 -88242 59962 -88208
rect 60000 -88242 60034 -88208
rect 60072 -88242 60106 -88208
rect 60144 -88242 60178 -88208
rect 60216 -88242 60250 -88208
rect 60288 -88242 60322 -88208
rect 60360 -88242 60394 -88208
rect 60432 -88242 60466 -88208
rect 60504 -88242 60538 -88208
rect 60576 -88242 60610 -88208
rect 60648 -88242 60682 -88208
rect 60720 -88242 60754 -88208
rect 60792 -88242 60826 -88208
rect 60864 -88242 60898 -88208
rect 60936 -88242 60970 -88208
rect 61008 -88242 61042 -88208
rect 61080 -88242 61114 -88208
rect 61152 -88242 61186 -88208
rect 61224 -88242 61258 -88208
rect 61296 -88242 61330 -88208
rect 61368 -88242 61402 -88208
rect 61440 -88242 61474 -88208
rect 61512 -88242 61546 -88208
rect 61584 -88242 61618 -88208
rect 61656 -88242 61690 -88208
rect 61728 -88242 61762 -88208
rect 61800 -88242 61834 -88208
rect 61872 -88242 61906 -88208
rect 61944 -88242 61978 -88208
rect 62016 -88242 62050 -88208
rect 62088 -88242 62122 -88208
rect 62160 -88242 62194 -88208
rect 62232 -88242 62266 -88208
rect 62304 -88242 62338 -88208
rect 62376 -88242 62410 -88208
rect 62448 -88242 62482 -88208
rect 62520 -88242 62554 -88208
rect 62592 -88242 62626 -88208
rect 62664 -88242 62698 -88208
rect 62736 -88242 62770 -88208
rect 62808 -88242 62842 -88208
rect 62880 -88242 62914 -88208
rect 62952 -88242 62986 -88208
rect 63024 -88242 63058 -88208
rect 63096 -88242 63130 -88208
rect 63168 -88242 63202 -88208
rect 63240 -88242 63274 -88208
rect 63312 -88242 63346 -88208
rect 63384 -88242 63418 -88208
rect 63456 -88242 63490 -88208
rect 63528 -88242 63562 -88208
rect 63600 -88242 63634 -88208
rect 63672 -88242 63706 -88208
rect 63744 -88242 63778 -88208
rect 63816 -88242 63850 -88208
rect 63888 -88242 63922 -88208
rect 63960 -88242 63994 -88208
rect 64032 -88242 64066 -88208
rect 64104 -88242 64138 -88208
rect 64176 -88242 64210 -88208
rect 64248 -88242 64282 -88208
<< metal1 >>
rect 52372 -69294 86359 -69270
rect 52372 -69390 68184 -69294
rect 52372 -69842 56256 -69390
rect 56130 -69858 56256 -69842
rect 64360 -69828 68184 -69390
rect 84246 -69828 86359 -69294
rect 64360 -69834 86359 -69828
rect 64360 -69858 86362 -69834
rect 56130 -69932 86362 -69858
rect 56294 -71294 56328 -69932
rect 56650 -71294 56684 -69932
rect 57006 -71294 57040 -69932
rect 57362 -71294 57396 -69932
rect 57718 -71292 57752 -69932
rect 58074 -71292 58108 -69932
rect 58432 -71292 58466 -69932
rect 58784 -71292 58818 -69932
rect 59142 -71292 59176 -69932
rect 59496 -71292 59530 -69932
rect 60786 -71288 60820 -69932
rect 60944 -71284 60954 -70132
rect 61012 -71284 61022 -70132
rect 61144 -71286 61178 -69932
rect 61300 -71286 61310 -70134
rect 61368 -71286 61378 -70134
rect 61500 -71288 61534 -69932
rect 61654 -71286 61664 -70134
rect 61722 -71286 61732 -70134
rect 61856 -71288 61890 -69932
rect 62012 -71280 62022 -70128
rect 62080 -71280 62090 -70128
rect 62210 -71284 62244 -69932
rect 62366 -71286 62376 -70134
rect 62434 -71286 62444 -70134
rect 62564 -71286 62598 -69932
rect 62720 -71284 62730 -70132
rect 62788 -71284 62798 -70132
rect 62922 -71284 62956 -69932
rect 63080 -71282 63090 -70130
rect 63148 -71282 63158 -70130
rect 63276 -71284 63310 -69932
rect 63436 -71284 63446 -70132
rect 63504 -71284 63514 -70132
rect 63634 -71280 63668 -69932
rect 63792 -71282 63802 -70130
rect 63860 -71282 63870 -70130
rect 63990 -71282 64024 -69932
rect 64150 -71282 64160 -70130
rect 64218 -71282 64228 -70130
rect 64348 -71278 64382 -69932
rect 68118 -71254 68128 -70112
rect 68182 -71254 68192 -70112
rect 68310 -71270 68320 -70128
rect 68374 -71270 68384 -70128
rect 68478 -71270 68488 -70128
rect 68542 -71270 68552 -70128
rect 68660 -71266 68670 -70124
rect 68724 -71266 68734 -70124
rect 68838 -71262 68848 -70120
rect 68902 -71262 68912 -70120
rect 69016 -71260 69026 -70118
rect 69080 -71260 69090 -70118
rect 69190 -71262 69200 -70120
rect 69254 -71262 69264 -70120
rect 69368 -71264 69378 -70122
rect 69432 -71264 69442 -70122
rect 69548 -71262 69558 -70120
rect 69612 -71262 69622 -70120
rect 69722 -71262 69732 -70120
rect 69786 -71262 69796 -70120
rect 69900 -71262 69910 -70120
rect 69964 -71262 69974 -70120
rect 70084 -71266 70094 -70124
rect 70148 -71266 70158 -70124
rect 70258 -71262 70268 -70120
rect 70322 -71262 70332 -70120
rect 70442 -71258 70452 -70116
rect 70506 -71258 70516 -70116
rect 70610 -71262 70620 -70120
rect 70674 -71262 70684 -70120
rect 70794 -71254 70804 -70112
rect 70858 -71254 70868 -70112
rect 70970 -71256 70980 -70114
rect 71034 -71256 71044 -70114
rect 71148 -71258 71158 -70116
rect 71212 -71258 71222 -70116
rect 71326 -71256 71336 -70114
rect 71390 -71256 71400 -70114
rect 71502 -71258 71512 -70116
rect 71566 -71258 71576 -70116
rect 71684 -71258 71694 -70116
rect 71748 -71258 71758 -70116
rect 71864 -71258 71874 -70116
rect 71928 -71258 71938 -70116
rect 72036 -71262 72046 -70120
rect 72100 -71262 72110 -70120
rect 72218 -71262 72228 -70120
rect 72282 -71262 72292 -70120
rect 72396 -71262 72406 -70120
rect 72460 -71262 72470 -70120
rect 72576 -71262 72586 -70120
rect 72640 -71262 72650 -70120
rect 72746 -71262 72756 -70120
rect 72810 -71262 72820 -70120
rect 72932 -71258 72942 -70116
rect 72996 -71258 73006 -70116
rect 73112 -71258 73122 -70116
rect 73176 -71258 73186 -70116
rect 73292 -71258 73302 -70116
rect 73356 -71258 73366 -70116
rect 73462 -71264 73472 -70122
rect 73526 -71264 73536 -70122
rect 73642 -71262 73652 -70120
rect 73706 -71262 73716 -70120
rect 73822 -71258 73832 -70116
rect 73886 -71258 73896 -70116
rect 73998 -71258 74008 -70116
rect 74062 -71258 74072 -70116
rect 74170 -71256 74180 -70114
rect 74234 -71256 74244 -70114
rect 74356 -71256 74366 -70114
rect 74420 -71256 74430 -70114
rect 74530 -71258 74540 -70116
rect 74594 -71258 74604 -70116
rect 74714 -71258 74724 -70116
rect 74778 -71258 74788 -70116
rect 74886 -71258 74896 -70116
rect 74950 -71258 74960 -70116
rect 75064 -71258 75074 -70116
rect 75128 -71258 75138 -70116
rect 75242 -71256 75252 -70114
rect 75306 -71256 75316 -70114
rect 75422 -71256 75432 -70114
rect 75486 -71256 75496 -70114
rect 75600 -71258 75610 -70116
rect 75664 -71258 75674 -70116
rect 75778 -71256 75788 -70114
rect 75842 -71256 75852 -70114
rect 75956 -71254 75966 -70112
rect 76020 -71254 76030 -70112
rect 76136 -71258 76146 -70116
rect 76200 -71258 76210 -70116
rect 76310 -71258 76320 -70116
rect 76374 -71258 76384 -70116
rect 76486 -71256 76496 -70114
rect 76550 -71256 76560 -70114
rect 76664 -71258 76674 -70116
rect 76728 -71258 76738 -70116
rect 76850 -71258 76860 -70116
rect 76914 -71258 76924 -70116
rect 77026 -71258 77036 -70116
rect 77090 -71258 77100 -70116
rect 77202 -71262 77212 -70120
rect 77266 -71262 77276 -70120
rect 77382 -71258 77392 -70116
rect 77446 -71258 77456 -70116
rect 77558 -71256 77568 -70114
rect 77622 -71256 77632 -70114
rect 77734 -71262 77744 -70120
rect 77798 -71262 77808 -70120
rect 77916 -71254 77926 -70112
rect 77980 -71254 77990 -70112
rect 78094 -71258 78104 -70116
rect 78158 -71258 78168 -70116
rect 78272 -71256 78282 -70114
rect 78336 -71256 78346 -70114
rect 78442 -71258 78452 -70116
rect 78506 -71258 78516 -70116
rect 78628 -71256 78638 -70114
rect 78692 -71256 78702 -70114
rect 78802 -71262 78812 -70120
rect 78866 -71262 78876 -70120
rect 78986 -71258 78996 -70116
rect 79050 -71258 79060 -70116
rect 79160 -71258 79170 -70116
rect 79224 -71258 79234 -70116
rect 79336 -71262 79346 -70120
rect 79400 -71262 79410 -70120
rect 79512 -71258 79522 -70116
rect 79576 -71258 79586 -70116
rect 79694 -71262 79704 -70120
rect 79758 -71262 79768 -70120
rect 79872 -71262 79882 -70120
rect 79936 -71262 79946 -70120
rect 80048 -71256 80058 -70114
rect 80112 -71256 80122 -70114
rect 80226 -71258 80236 -70116
rect 80290 -71258 80300 -70116
rect 80402 -71262 80412 -70120
rect 80466 -71262 80476 -70120
rect 80584 -71262 80594 -70120
rect 80648 -71262 80658 -70120
rect 80758 -71258 80768 -70116
rect 80822 -71258 80832 -70116
rect 80938 -71256 80948 -70114
rect 81002 -71256 81012 -70114
rect 81116 -71262 81126 -70120
rect 81180 -71262 81190 -70120
rect 81296 -71258 81306 -70116
rect 81360 -71258 81370 -70116
rect 81470 -71258 81480 -70116
rect 81534 -71258 81544 -70116
rect 81650 -71262 81660 -70120
rect 81714 -71262 81724 -70120
rect 81826 -71262 81836 -70120
rect 81890 -71262 81900 -70120
rect 82000 -71262 82010 -70120
rect 82064 -71262 82074 -70120
rect 82180 -71258 82190 -70116
rect 82244 -71258 82254 -70116
rect 82364 -71258 82374 -70116
rect 82428 -71258 82438 -70116
rect 82536 -71262 82546 -70120
rect 82600 -71262 82610 -70120
rect 82716 -71258 82726 -70116
rect 82780 -71258 82790 -70116
rect 82896 -71258 82906 -70116
rect 82960 -71258 82970 -70116
rect 83076 -71258 83086 -70116
rect 83140 -71258 83150 -70116
rect 83254 -71256 83264 -70114
rect 83318 -71256 83328 -70114
rect 83430 -71264 83440 -70122
rect 83494 -71264 83504 -70122
rect 83610 -71262 83620 -70120
rect 83674 -71262 83684 -70120
rect 83786 -71262 83796 -70120
rect 83850 -71262 83860 -70120
rect 83966 -71262 83976 -70120
rect 84030 -71262 84040 -70120
rect 84144 -71264 84154 -70122
rect 84208 -71264 84218 -70122
rect 68194 -71338 68204 -71328
rect 60836 -71343 60846 -71340
rect 60938 -71343 60948 -71340
rect 61192 -71343 61202 -71342
rect 61294 -71343 61304 -71342
rect 61548 -71343 61558 -71340
rect 61650 -71343 61660 -71340
rect 61726 -71343 61736 -71340
rect 61828 -71343 61838 -71340
rect 61906 -71343 61916 -71342
rect 62008 -71343 62018 -71342
rect 62080 -71343 62090 -71342
rect 62182 -71343 62192 -71342
rect 62438 -71343 62448 -71342
rect 62540 -71343 62550 -71342
rect 62800 -71343 62810 -71342
rect 62902 -71343 62912 -71342
rect 63328 -71343 63338 -71342
rect 63430 -71343 63440 -71342
rect 63684 -71343 63694 -71342
rect 63786 -71343 63796 -71342
rect 56320 -71484 56330 -71346
rect 59514 -71484 59524 -71346
rect 60824 -71482 60834 -71343
rect 64295 -71350 64305 -71343
rect 64320 -71406 64330 -71350
rect 64295 -71482 64305 -71406
rect 68190 -71482 68200 -71338
rect 68194 -71492 68204 -71482
rect 68302 -71492 68312 -71328
rect 68364 -71482 68374 -71338
rect 68470 -71482 68480 -71338
rect 68548 -71482 68558 -71338
rect 68654 -71482 68664 -71338
rect 68724 -71482 68734 -71338
rect 68830 -71482 68840 -71338
rect 68902 -71482 68912 -71338
rect 69008 -71482 69018 -71338
rect 69082 -71482 69092 -71338
rect 69188 -71482 69198 -71338
rect 69258 -71482 69268 -71338
rect 69364 -71482 69374 -71338
rect 69434 -71480 69444 -71336
rect 69540 -71480 69550 -71336
rect 69612 -71478 69622 -71334
rect 69718 -71478 69728 -71334
rect 69790 -71480 69800 -71336
rect 69896 -71480 69906 -71336
rect 69970 -71480 69980 -71336
rect 70076 -71480 70086 -71336
rect 70148 -71482 70158 -71338
rect 70254 -71482 70264 -71338
rect 70328 -71478 70338 -71334
rect 70434 -71478 70444 -71334
rect 70504 -71482 70514 -71338
rect 70610 -71482 70620 -71338
rect 70684 -71482 70694 -71338
rect 70790 -71482 70800 -71338
rect 70864 -71480 70874 -71336
rect 70970 -71480 70980 -71336
rect 71040 -71480 71050 -71336
rect 71146 -71480 71156 -71336
rect 71218 -71482 71228 -71338
rect 71324 -71482 71334 -71338
rect 71394 -71482 71404 -71338
rect 71500 -71482 71510 -71338
rect 71570 -71480 71580 -71336
rect 71676 -71480 71686 -71336
rect 71754 -71478 71764 -71334
rect 71860 -71478 71870 -71334
rect 71930 -71482 71940 -71338
rect 72036 -71482 72046 -71338
rect 72108 -71480 72118 -71336
rect 72214 -71480 72224 -71336
rect 72284 -71480 72294 -71336
rect 72390 -71480 72400 -71336
rect 72460 -71480 72470 -71336
rect 72566 -71480 72576 -71336
rect 72638 -71478 72648 -71334
rect 72744 -71478 72754 -71334
rect 72822 -71480 72832 -71336
rect 72928 -71480 72938 -71336
rect 72996 -71480 73006 -71336
rect 73102 -71480 73112 -71336
rect 73176 -71480 73186 -71336
rect 73282 -71480 73292 -71336
rect 73352 -71482 73362 -71338
rect 73458 -71482 73468 -71338
rect 73532 -71482 73542 -71338
rect 73638 -71482 73648 -71338
rect 73710 -71482 73720 -71338
rect 73816 -71482 73826 -71338
rect 73890 -71482 73900 -71338
rect 73996 -71482 74006 -71338
rect 74064 -71480 74074 -71336
rect 74170 -71480 74180 -71336
rect 74246 -71478 74256 -71334
rect 74352 -71478 74362 -71334
rect 74424 -71480 74434 -71336
rect 74530 -71480 74540 -71336
rect 74604 -71478 74614 -71334
rect 74710 -71478 74720 -71334
rect 74782 -71476 74792 -71332
rect 74888 -71476 74898 -71332
rect 74958 -71478 74968 -71334
rect 75064 -71478 75074 -71334
rect 75136 -71480 75146 -71336
rect 75242 -71480 75252 -71336
rect 75316 -71478 75326 -71334
rect 75422 -71478 75432 -71334
rect 75492 -71482 75502 -71338
rect 75598 -71482 75608 -71338
rect 75670 -71478 75680 -71334
rect 75776 -71478 75786 -71334
rect 75846 -71478 75856 -71334
rect 75952 -71478 75962 -71334
rect 76024 -71478 76034 -71334
rect 76130 -71478 76140 -71334
rect 76204 -71478 76214 -71334
rect 76310 -71478 76320 -71334
rect 76382 -71480 76392 -71336
rect 76488 -71480 76498 -71336
rect 76562 -71478 76572 -71334
rect 76668 -71478 76678 -71334
rect 76736 -71480 76746 -71336
rect 76842 -71480 76852 -71336
rect 76912 -71480 76922 -71336
rect 77018 -71480 77028 -71336
rect 77092 -71480 77102 -71336
rect 77198 -71480 77208 -71336
rect 77272 -71480 77282 -71336
rect 77378 -71480 77388 -71336
rect 77448 -71482 77458 -71338
rect 77554 -71482 77564 -71338
rect 77626 -71480 77636 -71336
rect 77732 -71480 77742 -71336
rect 77804 -71480 77814 -71336
rect 77910 -71480 77920 -71336
rect 77980 -71478 77990 -71334
rect 78086 -71478 78096 -71334
rect 78158 -71478 78168 -71334
rect 78264 -71478 78274 -71334
rect 78338 -71478 78348 -71334
rect 78444 -71478 78454 -71334
rect 78516 -71478 78526 -71334
rect 78622 -71478 78632 -71334
rect 78694 -71478 78704 -71334
rect 78800 -71478 78810 -71334
rect 78872 -71478 78882 -71334
rect 78978 -71478 78988 -71334
rect 79052 -71478 79062 -71334
rect 79158 -71478 79168 -71334
rect 79226 -71480 79236 -71336
rect 79332 -71480 79342 -71336
rect 79402 -71482 79412 -71338
rect 79508 -71482 79518 -71338
rect 79582 -71480 79592 -71336
rect 79688 -71480 79698 -71336
rect 79760 -71480 79770 -71336
rect 79866 -71480 79876 -71336
rect 79938 -71480 79948 -71336
rect 80044 -71480 80054 -71336
rect 80116 -71480 80126 -71336
rect 80222 -71480 80232 -71336
rect 80294 -71480 80304 -71336
rect 80400 -71480 80410 -71336
rect 80474 -71480 80484 -71336
rect 80580 -71480 80590 -71336
rect 80652 -71480 80662 -71336
rect 80758 -71480 80768 -71336
rect 80830 -71478 80840 -71334
rect 80936 -71478 80946 -71334
rect 81006 -71478 81016 -71334
rect 81112 -71478 81122 -71334
rect 81188 -71478 81198 -71334
rect 81294 -71478 81304 -71334
rect 81362 -71478 81372 -71334
rect 81468 -71478 81478 -71334
rect 81544 -71478 81554 -71334
rect 81650 -71478 81660 -71334
rect 81722 -71480 81732 -71336
rect 81828 -71480 81838 -71336
rect 81898 -71480 81908 -71336
rect 82004 -71480 82014 -71336
rect 82076 -71478 82086 -71334
rect 82182 -71478 82192 -71334
rect 82254 -71478 82264 -71334
rect 82360 -71478 82370 -71334
rect 82434 -71480 82444 -71336
rect 82540 -71480 82550 -71336
rect 82612 -71480 82622 -71336
rect 82718 -71480 82728 -71336
rect 82788 -71480 82798 -71336
rect 82894 -71480 82904 -71336
rect 82970 -71480 82980 -71336
rect 83076 -71480 83086 -71336
rect 83148 -71480 83158 -71336
rect 83254 -71480 83264 -71336
rect 83324 -71478 83334 -71334
rect 83430 -71478 83440 -71334
rect 83502 -71478 83512 -71334
rect 83608 -71478 83618 -71334
rect 83678 -71478 83688 -71334
rect 83784 -71478 83794 -71334
rect 83858 -71480 83868 -71336
rect 83964 -71480 83974 -71336
rect 84036 -71480 84046 -71336
rect 84142 -71480 84152 -71336
rect 68122 -72706 68132 -71562
rect 68190 -72706 68200 -71562
rect 68304 -72706 68314 -71562
rect 68372 -72706 68382 -71562
rect 68484 -72698 68494 -71554
rect 68552 -72698 68562 -71554
rect 68658 -72698 68668 -71554
rect 68726 -72698 68736 -71554
rect 68838 -72698 68848 -71554
rect 68906 -72698 68916 -71554
rect 69018 -72698 69028 -71554
rect 69086 -72698 69096 -71554
rect 69192 -72700 69202 -71556
rect 69260 -72700 69270 -71556
rect 69372 -72702 69382 -71558
rect 69440 -72702 69450 -71558
rect 69546 -72698 69556 -71554
rect 69614 -72698 69624 -71554
rect 69730 -72706 69740 -71562
rect 69798 -72706 69808 -71562
rect 69900 -72704 69910 -71560
rect 69968 -72704 69978 -71560
rect 70082 -72704 70092 -71560
rect 70150 -72704 70160 -71560
rect 70256 -72706 70266 -71562
rect 70324 -72706 70334 -71562
rect 70434 -72704 70444 -71560
rect 70502 -72704 70512 -71560
rect 70614 -72702 70624 -71558
rect 70682 -72702 70692 -71558
rect 70790 -72704 70800 -71560
rect 70858 -72704 70868 -71560
rect 70972 -72700 70982 -71556
rect 71040 -72700 71050 -71556
rect 71146 -72702 71156 -71558
rect 71214 -72702 71224 -71558
rect 71326 -72704 71336 -71560
rect 71394 -72704 71404 -71560
rect 71506 -72702 71516 -71558
rect 71574 -72702 71584 -71558
rect 71682 -72704 71692 -71560
rect 71750 -72704 71760 -71560
rect 71860 -72702 71870 -71558
rect 71928 -72702 71938 -71558
rect 72038 -72702 72048 -71558
rect 72106 -72702 72116 -71558
rect 72220 -72702 72230 -71558
rect 72288 -72702 72298 -71558
rect 72394 -72706 72404 -71562
rect 72462 -72706 72472 -71562
rect 72576 -72704 72586 -71560
rect 72644 -72704 72654 -71560
rect 72744 -72704 72754 -71560
rect 72812 -72704 72822 -71560
rect 72928 -72702 72938 -71558
rect 72996 -72702 73006 -71558
rect 73108 -72702 73118 -71558
rect 73176 -72702 73186 -71558
rect 73282 -72706 73292 -71562
rect 73350 -72706 73360 -71562
rect 73456 -72700 73466 -71556
rect 73524 -72700 73534 -71556
rect 73644 -72704 73654 -71560
rect 73712 -72704 73722 -71560
rect 73820 -72698 73830 -71554
rect 73888 -72698 73898 -71554
rect 74000 -72698 74010 -71554
rect 74068 -72698 74078 -71554
rect 74178 -72700 74188 -71556
rect 74246 -72700 74256 -71556
rect 74354 -72696 74364 -71552
rect 74422 -72696 74432 -71552
rect 74534 -72696 74544 -71552
rect 74602 -72696 74612 -71552
rect 74710 -72698 74720 -71554
rect 74778 -72698 74788 -71554
rect 74888 -72698 74898 -71554
rect 74956 -72698 74966 -71554
rect 75068 -72708 75078 -71564
rect 75136 -72708 75146 -71564
rect 75236 -72706 75246 -71562
rect 75304 -72706 75314 -71562
rect 75422 -72702 75432 -71558
rect 75490 -72702 75500 -71558
rect 75598 -72716 75608 -71572
rect 75666 -72716 75676 -71572
rect 75776 -72708 75786 -71564
rect 75844 -72708 75854 -71564
rect 75954 -72708 75964 -71564
rect 76022 -72708 76032 -71564
rect 76136 -72700 76146 -71556
rect 76204 -72700 76214 -71556
rect 76316 -72696 76326 -71552
rect 76384 -72696 76394 -71552
rect 76490 -72700 76500 -71556
rect 76558 -72700 76568 -71556
rect 76664 -72706 76674 -71562
rect 76732 -72706 76742 -71562
rect 76844 -72706 76854 -71562
rect 76912 -72706 76922 -71562
rect 77024 -72704 77034 -71560
rect 77092 -72704 77102 -71560
rect 77202 -72706 77212 -71562
rect 77270 -72706 77280 -71562
rect 77376 -72708 77386 -71564
rect 77444 -72708 77454 -71564
rect 77556 -72706 77566 -71562
rect 77624 -72706 77634 -71562
rect 77734 -72702 77744 -71558
rect 77802 -72702 77812 -71558
rect 77914 -72708 77924 -71564
rect 77982 -72708 77992 -71564
rect 78094 -72706 78104 -71562
rect 78162 -72706 78172 -71562
rect 78266 -72712 78276 -71568
rect 78334 -72712 78344 -71568
rect 78448 -72714 78458 -71570
rect 78516 -72714 78526 -71570
rect 78626 -72712 78636 -71568
rect 78694 -72712 78704 -71568
rect 78800 -72706 78810 -71562
rect 78868 -72706 78878 -71562
rect 78980 -72712 78990 -71568
rect 79048 -72712 79058 -71568
rect 79160 -72708 79170 -71564
rect 79228 -72708 79238 -71564
rect 79334 -72710 79344 -71566
rect 79402 -72710 79412 -71566
rect 79516 -72706 79526 -71562
rect 79584 -72706 79594 -71562
rect 79690 -72706 79700 -71562
rect 79758 -72706 79768 -71562
rect 79872 -72704 79882 -71560
rect 79940 -72704 79950 -71560
rect 80048 -72704 80058 -71560
rect 80116 -72704 80126 -71560
rect 80222 -72704 80232 -71560
rect 80290 -72704 80300 -71560
rect 80406 -72702 80416 -71558
rect 80474 -72702 80484 -71558
rect 80580 -72700 80590 -71556
rect 80648 -72700 80658 -71556
rect 80762 -72706 80772 -71562
rect 80830 -72706 80840 -71562
rect 80936 -72702 80946 -71558
rect 81004 -72702 81014 -71558
rect 81114 -72704 81124 -71560
rect 81182 -72704 81192 -71560
rect 81288 -72700 81298 -71556
rect 81356 -72700 81366 -71556
rect 81472 -72700 81482 -71556
rect 81540 -72700 81550 -71556
rect 81648 -72700 81658 -71556
rect 81716 -72700 81726 -71556
rect 81826 -72700 81836 -71556
rect 81894 -72700 81904 -71556
rect 82008 -72702 82018 -71558
rect 82076 -72702 82086 -71558
rect 82186 -72704 82196 -71560
rect 82254 -72704 82264 -71560
rect 82360 -72706 82370 -71562
rect 82428 -72706 82438 -71562
rect 82546 -72702 82556 -71558
rect 82614 -72702 82624 -71558
rect 82714 -72704 82724 -71560
rect 82782 -72704 82792 -71560
rect 82898 -72698 82908 -71554
rect 82966 -72698 82976 -71554
rect 83070 -72698 83080 -71554
rect 83138 -72698 83148 -71554
rect 83252 -72698 83262 -71554
rect 83320 -72698 83330 -71554
rect 83434 -72704 83444 -71560
rect 83502 -72704 83512 -71560
rect 83612 -72706 83622 -71562
rect 83680 -72706 83690 -71562
rect 83786 -72706 83796 -71562
rect 83854 -72706 83864 -71562
rect 83968 -72700 83978 -71556
rect 84036 -72700 84046 -71556
rect 84138 -72710 84148 -71566
rect 84206 -72710 84216 -71566
rect 84400 -72866 86362 -69932
rect 55932 -73126 56350 -72922
rect 56304 -74544 56314 -73398
rect 56368 -74544 56378 -73398
rect 56480 -74542 56490 -73396
rect 56544 -74542 56554 -73396
rect 56658 -74546 56668 -73400
rect 56722 -74546 56732 -73400
rect 56842 -74542 56852 -73396
rect 56906 -74542 56916 -73396
rect 57016 -74550 57026 -73404
rect 57080 -74550 57090 -73404
rect 57192 -74554 57202 -73408
rect 57256 -74554 57266 -73408
rect 57372 -74550 57382 -73404
rect 57436 -74550 57446 -73404
rect 57548 -74546 57558 -73400
rect 57612 -74546 57622 -73400
rect 57730 -74546 57740 -73400
rect 57794 -74546 57804 -73400
rect 57906 -74550 57916 -73404
rect 57970 -74550 57980 -73404
rect 58084 -74550 58094 -73404
rect 58148 -74550 58158 -73404
rect 58266 -74554 58276 -73408
rect 58330 -74554 58340 -73408
rect 58440 -74550 58450 -73404
rect 58504 -74550 58514 -73404
rect 58620 -74548 58630 -73402
rect 58684 -74548 58694 -73402
rect 58796 -74548 58806 -73402
rect 58860 -74548 58870 -73402
rect 58976 -74546 58986 -73400
rect 59040 -74546 59050 -73400
rect 59156 -74546 59166 -73400
rect 59220 -74546 59230 -73400
rect 59334 -74546 59344 -73400
rect 59398 -74546 59408 -73400
rect 59512 -74542 59522 -73396
rect 59576 -74542 59586 -73396
rect 59688 -74546 59698 -73400
rect 59752 -74546 59762 -73400
rect 59866 -74550 59876 -73404
rect 59930 -74550 59940 -73404
rect 60044 -74550 60054 -73404
rect 60108 -74550 60118 -73404
rect 60218 -74550 60228 -73404
rect 60282 -74550 60292 -73404
rect 60396 -74554 60406 -73408
rect 60460 -74554 60470 -73408
rect 60578 -74554 60588 -73408
rect 60642 -74554 60652 -73408
rect 60758 -74546 60768 -73400
rect 60822 -74546 60832 -73400
rect 60934 -74550 60944 -73404
rect 60998 -74550 61008 -73404
rect 61112 -74550 61122 -73404
rect 61176 -74550 61186 -73404
rect 61288 -74554 61298 -73408
rect 61352 -74554 61362 -73408
rect 61468 -74548 61478 -73402
rect 61532 -74548 61542 -73402
rect 61646 -74546 61656 -73400
rect 61710 -74546 61720 -73400
rect 61818 -74550 61828 -73404
rect 61882 -74550 61892 -73404
rect 61998 -74550 62008 -73404
rect 62062 -74550 62072 -73404
rect 62178 -74550 62188 -73404
rect 62242 -74550 62252 -73404
rect 62358 -74550 62368 -73404
rect 62422 -74550 62432 -73404
rect 62536 -74548 62546 -73402
rect 62600 -74548 62610 -73402
rect 62710 -74544 62720 -73398
rect 62774 -74544 62784 -73398
rect 62888 -74550 62898 -73404
rect 62952 -74550 62962 -73404
rect 63070 -74548 63080 -73402
rect 63134 -74548 63144 -73402
rect 63246 -74544 63256 -73398
rect 63310 -74544 63320 -73398
rect 63422 -74548 63432 -73402
rect 63486 -74548 63496 -73402
rect 63602 -74546 63612 -73400
rect 63666 -74546 63676 -73400
rect 63780 -74546 63790 -73400
rect 63844 -74546 63854 -73400
rect 63958 -74544 63968 -73398
rect 64022 -74544 64032 -73398
rect 64136 -74542 64146 -73396
rect 64200 -74542 64210 -73396
rect 64312 -74546 64322 -73400
rect 64376 -74546 64386 -73400
rect 56354 -74792 56364 -74636
rect 56470 -74792 56480 -74636
rect 56536 -74798 56546 -74642
rect 56652 -74798 56662 -74642
rect 56718 -74794 56728 -74638
rect 56834 -74794 56844 -74638
rect 56898 -74794 56908 -74638
rect 57014 -74794 57024 -74638
rect 57076 -74792 57086 -74636
rect 57192 -74792 57202 -74636
rect 57252 -74792 57262 -74636
rect 57368 -74792 57378 -74636
rect 57436 -74794 57446 -74638
rect 57552 -74794 57562 -74638
rect 57610 -74794 57620 -74638
rect 57726 -74794 57736 -74638
rect 57784 -74794 57794 -74638
rect 57900 -74794 57910 -74638
rect 57966 -74798 57976 -74642
rect 58082 -74798 58092 -74642
rect 58140 -74794 58150 -74638
rect 58256 -74794 58266 -74638
rect 58318 -74794 58328 -74638
rect 58434 -74794 58444 -74638
rect 58498 -74794 58508 -74638
rect 58614 -74794 58624 -74638
rect 58668 -74794 58678 -74638
rect 58784 -74794 58794 -74638
rect 58848 -74794 58858 -74638
rect 58964 -74794 58974 -74638
rect 59032 -74794 59042 -74638
rect 59148 -74794 59158 -74638
rect 59206 -74794 59216 -74638
rect 59322 -74794 59332 -74638
rect 59380 -74792 59390 -74636
rect 59496 -74792 59506 -74636
rect 59558 -74788 59568 -74632
rect 59674 -74788 59684 -74632
rect 59740 -74798 59750 -74642
rect 59856 -74798 59866 -74642
rect 59916 -74794 59926 -74638
rect 60032 -74794 60042 -74638
rect 60096 -74794 60106 -74638
rect 60212 -74794 60222 -74638
rect 60268 -74794 60278 -74638
rect 60384 -74794 60394 -74638
rect 60452 -74798 60462 -74642
rect 60568 -74798 60578 -74642
rect 60626 -74794 60636 -74638
rect 60742 -74794 60752 -74638
rect 60806 -74798 60816 -74642
rect 60922 -74798 60932 -74642
rect 60982 -74798 60992 -74642
rect 61098 -74798 61108 -74642
rect 61158 -74794 61168 -74638
rect 61274 -74794 61284 -74638
rect 61338 -74798 61348 -74642
rect 61454 -74798 61464 -74642
rect 61518 -74794 61528 -74638
rect 61634 -74794 61644 -74638
rect 61696 -74802 61706 -74646
rect 61812 -74802 61822 -74646
rect 61876 -74794 61886 -74638
rect 61992 -74794 62002 -74638
rect 62052 -74798 62062 -74642
rect 62168 -74798 62178 -74642
rect 62230 -74788 62240 -74632
rect 62346 -74788 62356 -74632
rect 62408 -74794 62418 -74638
rect 62524 -74794 62534 -74638
rect 62586 -74794 62596 -74638
rect 62702 -74794 62712 -74638
rect 62766 -74798 62776 -74642
rect 62882 -74798 62892 -74642
rect 62946 -74798 62956 -74642
rect 63062 -74798 63072 -74642
rect 63120 -74794 63130 -74638
rect 63236 -74794 63246 -74638
rect 63304 -74798 63314 -74642
rect 63420 -74798 63430 -74642
rect 63472 -74798 63482 -74642
rect 63588 -74798 63598 -74642
rect 63650 -74804 63660 -74648
rect 63766 -74804 63776 -74648
rect 63838 -74792 63848 -74636
rect 63954 -74792 63964 -74636
rect 64010 -74794 64020 -74638
rect 64126 -74794 64136 -74638
rect 64190 -74792 64200 -74636
rect 64306 -74792 64316 -74636
rect 56288 -76006 56298 -74860
rect 56352 -76006 56362 -74860
rect 56464 -76004 56474 -74858
rect 56528 -76004 56538 -74858
rect 56642 -76008 56652 -74862
rect 56706 -76008 56716 -74862
rect 56826 -76004 56836 -74858
rect 56890 -76004 56900 -74858
rect 57000 -76012 57010 -74866
rect 57064 -76012 57074 -74866
rect 57176 -76016 57186 -74870
rect 57240 -76016 57250 -74870
rect 57356 -76012 57366 -74866
rect 57420 -76012 57430 -74866
rect 57532 -76008 57542 -74862
rect 57596 -76008 57606 -74862
rect 57714 -76008 57724 -74862
rect 57778 -76008 57788 -74862
rect 57890 -76012 57900 -74866
rect 57954 -76012 57964 -74866
rect 58068 -76012 58078 -74866
rect 58132 -76012 58142 -74866
rect 58250 -76016 58260 -74870
rect 58314 -76016 58324 -74870
rect 58424 -76012 58434 -74866
rect 58488 -76012 58498 -74866
rect 58604 -76010 58614 -74864
rect 58668 -76010 58678 -74864
rect 58780 -76010 58790 -74864
rect 58844 -76010 58854 -74864
rect 58960 -76008 58970 -74862
rect 59024 -76008 59034 -74862
rect 59140 -76008 59150 -74862
rect 59204 -76008 59214 -74862
rect 59318 -76008 59328 -74862
rect 59382 -76008 59392 -74862
rect 59496 -76004 59506 -74858
rect 59560 -76004 59570 -74858
rect 59672 -76008 59682 -74862
rect 59736 -76008 59746 -74862
rect 59850 -76012 59860 -74866
rect 59914 -76012 59924 -74866
rect 60028 -76012 60038 -74866
rect 60092 -76012 60102 -74866
rect 60202 -76012 60212 -74866
rect 60266 -76012 60276 -74866
rect 60380 -76016 60390 -74870
rect 60444 -76016 60454 -74870
rect 60562 -76016 60572 -74870
rect 60626 -76016 60636 -74870
rect 60742 -76008 60752 -74862
rect 60806 -76008 60816 -74862
rect 60918 -76012 60928 -74866
rect 60982 -76012 60992 -74866
rect 61096 -76012 61106 -74866
rect 61160 -76012 61170 -74866
rect 61272 -76016 61282 -74870
rect 61336 -76016 61346 -74870
rect 61452 -76010 61462 -74864
rect 61516 -76010 61526 -74864
rect 61630 -76008 61640 -74862
rect 61694 -76008 61704 -74862
rect 61802 -76012 61812 -74866
rect 61866 -76012 61876 -74866
rect 61982 -76012 61992 -74866
rect 62046 -76012 62056 -74866
rect 62162 -76012 62172 -74866
rect 62226 -76012 62236 -74866
rect 62342 -76012 62352 -74866
rect 62406 -76012 62416 -74866
rect 62520 -76010 62530 -74864
rect 62584 -76010 62594 -74864
rect 62694 -76006 62704 -74860
rect 62758 -76006 62768 -74860
rect 62872 -76012 62882 -74866
rect 62936 -76012 62946 -74866
rect 63054 -76010 63064 -74864
rect 63118 -76010 63128 -74864
rect 63230 -76006 63240 -74860
rect 63294 -76006 63304 -74860
rect 63406 -76010 63416 -74864
rect 63470 -76010 63480 -74864
rect 63586 -76008 63596 -74862
rect 63650 -76008 63660 -74862
rect 63764 -76008 63774 -74862
rect 63828 -76008 63838 -74862
rect 63942 -76006 63952 -74860
rect 64006 -76006 64016 -74860
rect 64120 -76004 64130 -74858
rect 64184 -76004 64194 -74858
rect 64296 -76008 64306 -74862
rect 64360 -76008 64370 -74862
rect 56032 -76728 56326 -76506
rect 56294 -78394 56304 -77248
rect 56358 -78394 56368 -77248
rect 56470 -78392 56480 -77246
rect 56534 -78392 56544 -77246
rect 56648 -78396 56658 -77250
rect 56712 -78396 56722 -77250
rect 56832 -78392 56842 -77246
rect 56896 -78392 56906 -77246
rect 57006 -78400 57016 -77254
rect 57070 -78400 57080 -77254
rect 57182 -78404 57192 -77258
rect 57246 -78404 57256 -77258
rect 57362 -78400 57372 -77254
rect 57426 -78400 57436 -77254
rect 57538 -78396 57548 -77250
rect 57602 -78396 57612 -77250
rect 57720 -78396 57730 -77250
rect 57784 -78396 57794 -77250
rect 57896 -78400 57906 -77254
rect 57960 -78400 57970 -77254
rect 58074 -78400 58084 -77254
rect 58138 -78400 58148 -77254
rect 58256 -78404 58266 -77258
rect 58320 -78404 58330 -77258
rect 58430 -78400 58440 -77254
rect 58494 -78400 58504 -77254
rect 58610 -78398 58620 -77252
rect 58674 -78398 58684 -77252
rect 58786 -78398 58796 -77252
rect 58850 -78398 58860 -77252
rect 58966 -78396 58976 -77250
rect 59030 -78396 59040 -77250
rect 59146 -78396 59156 -77250
rect 59210 -78396 59220 -77250
rect 59324 -78396 59334 -77250
rect 59388 -78396 59398 -77250
rect 59502 -78392 59512 -77246
rect 59566 -78392 59576 -77246
rect 59678 -78396 59688 -77250
rect 59742 -78396 59752 -77250
rect 59856 -78400 59866 -77254
rect 59920 -78400 59930 -77254
rect 60034 -78400 60044 -77254
rect 60098 -78400 60108 -77254
rect 60208 -78400 60218 -77254
rect 60272 -78400 60282 -77254
rect 60386 -78404 60396 -77258
rect 60450 -78404 60460 -77258
rect 60568 -78404 60578 -77258
rect 60632 -78404 60642 -77258
rect 60748 -78396 60758 -77250
rect 60812 -78396 60822 -77250
rect 60924 -78400 60934 -77254
rect 60988 -78400 60998 -77254
rect 61102 -78400 61112 -77254
rect 61166 -78400 61176 -77254
rect 61278 -78404 61288 -77258
rect 61342 -78404 61352 -77258
rect 61458 -78398 61468 -77252
rect 61522 -78398 61532 -77252
rect 61636 -78396 61646 -77250
rect 61700 -78396 61710 -77250
rect 61808 -78400 61818 -77254
rect 61872 -78400 61882 -77254
rect 61988 -78400 61998 -77254
rect 62052 -78400 62062 -77254
rect 62168 -78400 62178 -77254
rect 62232 -78400 62242 -77254
rect 62348 -78400 62358 -77254
rect 62412 -78400 62422 -77254
rect 62526 -78398 62536 -77252
rect 62590 -78398 62600 -77252
rect 62700 -78394 62710 -77248
rect 62764 -78394 62774 -77248
rect 62878 -78400 62888 -77254
rect 62942 -78400 62952 -77254
rect 63060 -78398 63070 -77252
rect 63124 -78398 63134 -77252
rect 63236 -78394 63246 -77248
rect 63300 -78394 63310 -77248
rect 63412 -78398 63422 -77252
rect 63476 -78398 63486 -77252
rect 63592 -78396 63602 -77250
rect 63656 -78396 63666 -77250
rect 63770 -78396 63780 -77250
rect 63834 -78396 63844 -77250
rect 63948 -78394 63958 -77248
rect 64012 -78394 64022 -77248
rect 64126 -78392 64136 -77246
rect 64190 -78392 64200 -77246
rect 64302 -78396 64312 -77250
rect 64366 -78396 64376 -77250
rect 56344 -78642 56354 -78486
rect 56460 -78642 56470 -78486
rect 56526 -78648 56536 -78492
rect 56642 -78648 56652 -78492
rect 56708 -78644 56718 -78488
rect 56824 -78644 56834 -78488
rect 56888 -78644 56898 -78488
rect 57004 -78644 57014 -78488
rect 57066 -78642 57076 -78486
rect 57182 -78642 57192 -78486
rect 57242 -78642 57252 -78486
rect 57358 -78642 57368 -78486
rect 57426 -78644 57436 -78488
rect 57542 -78644 57552 -78488
rect 57600 -78644 57610 -78488
rect 57716 -78644 57726 -78488
rect 57774 -78644 57784 -78488
rect 57890 -78644 57900 -78488
rect 57956 -78648 57966 -78492
rect 58072 -78648 58082 -78492
rect 58130 -78644 58140 -78488
rect 58246 -78644 58256 -78488
rect 58308 -78644 58318 -78488
rect 58424 -78644 58434 -78488
rect 58488 -78644 58498 -78488
rect 58604 -78644 58614 -78488
rect 58658 -78644 58668 -78488
rect 58774 -78644 58784 -78488
rect 58838 -78644 58848 -78488
rect 58954 -78644 58964 -78488
rect 59022 -78644 59032 -78488
rect 59138 -78644 59148 -78488
rect 59196 -78644 59206 -78488
rect 59312 -78644 59322 -78488
rect 59370 -78642 59380 -78486
rect 59486 -78642 59496 -78486
rect 59548 -78638 59558 -78482
rect 59664 -78638 59674 -78482
rect 59730 -78648 59740 -78492
rect 59846 -78648 59856 -78492
rect 59906 -78644 59916 -78488
rect 60022 -78644 60032 -78488
rect 60086 -78644 60096 -78488
rect 60202 -78644 60212 -78488
rect 60258 -78644 60268 -78488
rect 60374 -78644 60384 -78488
rect 60442 -78648 60452 -78492
rect 60558 -78648 60568 -78492
rect 60616 -78644 60626 -78488
rect 60732 -78644 60742 -78488
rect 60796 -78648 60806 -78492
rect 60912 -78648 60922 -78492
rect 60972 -78648 60982 -78492
rect 61088 -78648 61098 -78492
rect 61148 -78644 61158 -78488
rect 61264 -78644 61274 -78488
rect 61328 -78648 61338 -78492
rect 61444 -78648 61454 -78492
rect 61508 -78644 61518 -78488
rect 61624 -78644 61634 -78488
rect 61686 -78652 61696 -78496
rect 61802 -78652 61812 -78496
rect 61866 -78644 61876 -78488
rect 61982 -78644 61992 -78488
rect 62042 -78648 62052 -78492
rect 62158 -78648 62168 -78492
rect 62220 -78638 62230 -78482
rect 62336 -78638 62346 -78482
rect 62398 -78644 62408 -78488
rect 62514 -78644 62524 -78488
rect 62576 -78644 62586 -78488
rect 62692 -78644 62702 -78488
rect 62756 -78648 62766 -78492
rect 62872 -78648 62882 -78492
rect 62936 -78648 62946 -78492
rect 63052 -78648 63062 -78492
rect 63110 -78644 63120 -78488
rect 63226 -78644 63236 -78488
rect 63294 -78648 63304 -78492
rect 63410 -78648 63420 -78492
rect 63462 -78648 63472 -78492
rect 63578 -78648 63588 -78492
rect 63640 -78654 63650 -78498
rect 63756 -78654 63766 -78498
rect 63828 -78642 63838 -78486
rect 63944 -78642 63954 -78486
rect 64000 -78644 64010 -78488
rect 64116 -78644 64126 -78488
rect 64180 -78642 64190 -78486
rect 64296 -78642 64306 -78486
rect 56278 -79856 56288 -78710
rect 56342 -79856 56352 -78710
rect 56454 -79854 56464 -78708
rect 56518 -79854 56528 -78708
rect 56632 -79858 56642 -78712
rect 56696 -79858 56706 -78712
rect 56816 -79854 56826 -78708
rect 56880 -79854 56890 -78708
rect 56990 -79862 57000 -78716
rect 57054 -79862 57064 -78716
rect 57166 -79866 57176 -78720
rect 57230 -79866 57240 -78720
rect 57346 -79862 57356 -78716
rect 57410 -79862 57420 -78716
rect 57522 -79858 57532 -78712
rect 57586 -79858 57596 -78712
rect 57704 -79858 57714 -78712
rect 57768 -79858 57778 -78712
rect 57880 -79862 57890 -78716
rect 57944 -79862 57954 -78716
rect 58058 -79862 58068 -78716
rect 58122 -79862 58132 -78716
rect 58240 -79866 58250 -78720
rect 58304 -79866 58314 -78720
rect 58414 -79862 58424 -78716
rect 58478 -79862 58488 -78716
rect 58594 -79860 58604 -78714
rect 58658 -79860 58668 -78714
rect 58770 -79860 58780 -78714
rect 58834 -79860 58844 -78714
rect 58950 -79858 58960 -78712
rect 59014 -79858 59024 -78712
rect 59130 -79858 59140 -78712
rect 59194 -79858 59204 -78712
rect 59308 -79858 59318 -78712
rect 59372 -79858 59382 -78712
rect 59486 -79854 59496 -78708
rect 59550 -79854 59560 -78708
rect 59662 -79858 59672 -78712
rect 59726 -79858 59736 -78712
rect 59840 -79862 59850 -78716
rect 59904 -79862 59914 -78716
rect 60018 -79862 60028 -78716
rect 60082 -79862 60092 -78716
rect 60192 -79862 60202 -78716
rect 60256 -79862 60266 -78716
rect 60370 -79866 60380 -78720
rect 60434 -79866 60444 -78720
rect 60552 -79866 60562 -78720
rect 60616 -79866 60626 -78720
rect 60732 -79858 60742 -78712
rect 60796 -79858 60806 -78712
rect 60908 -79862 60918 -78716
rect 60972 -79862 60982 -78716
rect 61086 -79862 61096 -78716
rect 61150 -79862 61160 -78716
rect 61262 -79866 61272 -78720
rect 61326 -79866 61336 -78720
rect 61442 -79860 61452 -78714
rect 61506 -79860 61516 -78714
rect 61620 -79858 61630 -78712
rect 61684 -79858 61694 -78712
rect 61792 -79862 61802 -78716
rect 61856 -79862 61866 -78716
rect 61972 -79862 61982 -78716
rect 62036 -79862 62046 -78716
rect 62152 -79862 62162 -78716
rect 62216 -79862 62226 -78716
rect 62332 -79862 62342 -78716
rect 62396 -79862 62406 -78716
rect 62510 -79860 62520 -78714
rect 62574 -79860 62584 -78714
rect 62684 -79856 62694 -78710
rect 62748 -79856 62758 -78710
rect 62862 -79862 62872 -78716
rect 62926 -79862 62936 -78716
rect 63044 -79860 63054 -78714
rect 63108 -79860 63118 -78714
rect 63220 -79856 63230 -78710
rect 63284 -79856 63294 -78710
rect 63396 -79860 63406 -78714
rect 63460 -79860 63470 -78714
rect 63576 -79858 63586 -78712
rect 63640 -79858 63650 -78712
rect 63754 -79858 63764 -78712
rect 63818 -79858 63828 -78712
rect 63932 -79856 63942 -78710
rect 63996 -79856 64006 -78710
rect 64110 -79854 64120 -78708
rect 64174 -79854 64184 -78708
rect 64286 -79858 64296 -78712
rect 64350 -79858 64360 -78712
rect 56028 -80712 56322 -80490
rect 56304 -82360 56314 -81214
rect 56368 -82360 56378 -81214
rect 56480 -82358 56490 -81212
rect 56544 -82358 56554 -81212
rect 56658 -82362 56668 -81216
rect 56722 -82362 56732 -81216
rect 56842 -82358 56852 -81212
rect 56906 -82358 56916 -81212
rect 57016 -82366 57026 -81220
rect 57080 -82366 57090 -81220
rect 57192 -82370 57202 -81224
rect 57256 -82370 57266 -81224
rect 57372 -82366 57382 -81220
rect 57436 -82366 57446 -81220
rect 57548 -82362 57558 -81216
rect 57612 -82362 57622 -81216
rect 57730 -82362 57740 -81216
rect 57794 -82362 57804 -81216
rect 57906 -82366 57916 -81220
rect 57970 -82366 57980 -81220
rect 58084 -82366 58094 -81220
rect 58148 -82366 58158 -81220
rect 58266 -82370 58276 -81224
rect 58330 -82370 58340 -81224
rect 58440 -82366 58450 -81220
rect 58504 -82366 58514 -81220
rect 58620 -82364 58630 -81218
rect 58684 -82364 58694 -81218
rect 58796 -82364 58806 -81218
rect 58860 -82364 58870 -81218
rect 58976 -82362 58986 -81216
rect 59040 -82362 59050 -81216
rect 59156 -82362 59166 -81216
rect 59220 -82362 59230 -81216
rect 59334 -82362 59344 -81216
rect 59398 -82362 59408 -81216
rect 59512 -82358 59522 -81212
rect 59576 -82358 59586 -81212
rect 59688 -82362 59698 -81216
rect 59752 -82362 59762 -81216
rect 59866 -82366 59876 -81220
rect 59930 -82366 59940 -81220
rect 60044 -82366 60054 -81220
rect 60108 -82366 60118 -81220
rect 60218 -82366 60228 -81220
rect 60282 -82366 60292 -81220
rect 60396 -82370 60406 -81224
rect 60460 -82370 60470 -81224
rect 60578 -82370 60588 -81224
rect 60642 -82370 60652 -81224
rect 60758 -82362 60768 -81216
rect 60822 -82362 60832 -81216
rect 60934 -82366 60944 -81220
rect 60998 -82366 61008 -81220
rect 61112 -82366 61122 -81220
rect 61176 -82366 61186 -81220
rect 61288 -82370 61298 -81224
rect 61352 -82370 61362 -81224
rect 61468 -82364 61478 -81218
rect 61532 -82364 61542 -81218
rect 61646 -82362 61656 -81216
rect 61710 -82362 61720 -81216
rect 61818 -82366 61828 -81220
rect 61882 -82366 61892 -81220
rect 61998 -82366 62008 -81220
rect 62062 -82366 62072 -81220
rect 62178 -82366 62188 -81220
rect 62242 -82366 62252 -81220
rect 62358 -82366 62368 -81220
rect 62422 -82366 62432 -81220
rect 62536 -82364 62546 -81218
rect 62600 -82364 62610 -81218
rect 62710 -82360 62720 -81214
rect 62774 -82360 62784 -81214
rect 62888 -82366 62898 -81220
rect 62952 -82366 62962 -81220
rect 63070 -82364 63080 -81218
rect 63134 -82364 63144 -81218
rect 63246 -82360 63256 -81214
rect 63310 -82360 63320 -81214
rect 63422 -82364 63432 -81218
rect 63486 -82364 63496 -81218
rect 63602 -82362 63612 -81216
rect 63666 -82362 63676 -81216
rect 63780 -82362 63790 -81216
rect 63844 -82362 63854 -81216
rect 63958 -82360 63968 -81214
rect 64022 -82360 64032 -81214
rect 64136 -82358 64146 -81212
rect 64200 -82358 64210 -81212
rect 64312 -82362 64322 -81216
rect 64376 -82362 64386 -81216
rect 56354 -82608 56364 -82452
rect 56470 -82608 56480 -82452
rect 56536 -82614 56546 -82458
rect 56652 -82614 56662 -82458
rect 56718 -82610 56728 -82454
rect 56834 -82610 56844 -82454
rect 56898 -82610 56908 -82454
rect 57014 -82610 57024 -82454
rect 57076 -82608 57086 -82452
rect 57192 -82608 57202 -82452
rect 57252 -82608 57262 -82452
rect 57368 -82608 57378 -82452
rect 57436 -82610 57446 -82454
rect 57552 -82610 57562 -82454
rect 57610 -82610 57620 -82454
rect 57726 -82610 57736 -82454
rect 57784 -82610 57794 -82454
rect 57900 -82610 57910 -82454
rect 57966 -82614 57976 -82458
rect 58082 -82614 58092 -82458
rect 58140 -82610 58150 -82454
rect 58256 -82610 58266 -82454
rect 58318 -82610 58328 -82454
rect 58434 -82610 58444 -82454
rect 58498 -82610 58508 -82454
rect 58614 -82610 58624 -82454
rect 58668 -82610 58678 -82454
rect 58784 -82610 58794 -82454
rect 58848 -82610 58858 -82454
rect 58964 -82610 58974 -82454
rect 59032 -82610 59042 -82454
rect 59148 -82610 59158 -82454
rect 59206 -82610 59216 -82454
rect 59322 -82610 59332 -82454
rect 59380 -82608 59390 -82452
rect 59496 -82608 59506 -82452
rect 59558 -82604 59568 -82448
rect 59674 -82604 59684 -82448
rect 59740 -82614 59750 -82458
rect 59856 -82614 59866 -82458
rect 59916 -82610 59926 -82454
rect 60032 -82610 60042 -82454
rect 60096 -82610 60106 -82454
rect 60212 -82610 60222 -82454
rect 60268 -82610 60278 -82454
rect 60384 -82610 60394 -82454
rect 60452 -82614 60462 -82458
rect 60568 -82614 60578 -82458
rect 60626 -82610 60636 -82454
rect 60742 -82610 60752 -82454
rect 60806 -82614 60816 -82458
rect 60922 -82614 60932 -82458
rect 60982 -82614 60992 -82458
rect 61098 -82614 61108 -82458
rect 61158 -82610 61168 -82454
rect 61274 -82610 61284 -82454
rect 61338 -82614 61348 -82458
rect 61454 -82614 61464 -82458
rect 61518 -82610 61528 -82454
rect 61634 -82610 61644 -82454
rect 61696 -82618 61706 -82462
rect 61812 -82618 61822 -82462
rect 61876 -82610 61886 -82454
rect 61992 -82610 62002 -82454
rect 62052 -82614 62062 -82458
rect 62168 -82614 62178 -82458
rect 62230 -82604 62240 -82448
rect 62346 -82604 62356 -82448
rect 62408 -82610 62418 -82454
rect 62524 -82610 62534 -82454
rect 62586 -82610 62596 -82454
rect 62702 -82610 62712 -82454
rect 62766 -82614 62776 -82458
rect 62882 -82614 62892 -82458
rect 62946 -82614 62956 -82458
rect 63062 -82614 63072 -82458
rect 63120 -82610 63130 -82454
rect 63236 -82610 63246 -82454
rect 63304 -82614 63314 -82458
rect 63420 -82614 63430 -82458
rect 63472 -82614 63482 -82458
rect 63588 -82614 63598 -82458
rect 63650 -82620 63660 -82464
rect 63766 -82620 63776 -82464
rect 63838 -82608 63848 -82452
rect 63954 -82608 63964 -82452
rect 64010 -82610 64020 -82454
rect 64126 -82610 64136 -82454
rect 64190 -82608 64200 -82452
rect 64306 -82608 64316 -82452
rect 56288 -83822 56298 -82676
rect 56352 -83822 56362 -82676
rect 56464 -83820 56474 -82674
rect 56528 -83820 56538 -82674
rect 56642 -83824 56652 -82678
rect 56706 -83824 56716 -82678
rect 56826 -83820 56836 -82674
rect 56890 -83820 56900 -82674
rect 57000 -83828 57010 -82682
rect 57064 -83828 57074 -82682
rect 57176 -83832 57186 -82686
rect 57240 -83832 57250 -82686
rect 57356 -83828 57366 -82682
rect 57420 -83828 57430 -82682
rect 57532 -83824 57542 -82678
rect 57596 -83824 57606 -82678
rect 57714 -83824 57724 -82678
rect 57778 -83824 57788 -82678
rect 57890 -83828 57900 -82682
rect 57954 -83828 57964 -82682
rect 58068 -83828 58078 -82682
rect 58132 -83828 58142 -82682
rect 58250 -83832 58260 -82686
rect 58314 -83832 58324 -82686
rect 58424 -83828 58434 -82682
rect 58488 -83828 58498 -82682
rect 58604 -83826 58614 -82680
rect 58668 -83826 58678 -82680
rect 58780 -83826 58790 -82680
rect 58844 -83826 58854 -82680
rect 58960 -83824 58970 -82678
rect 59024 -83824 59034 -82678
rect 59140 -83824 59150 -82678
rect 59204 -83824 59214 -82678
rect 59318 -83824 59328 -82678
rect 59382 -83824 59392 -82678
rect 59496 -83820 59506 -82674
rect 59560 -83820 59570 -82674
rect 59672 -83824 59682 -82678
rect 59736 -83824 59746 -82678
rect 59850 -83828 59860 -82682
rect 59914 -83828 59924 -82682
rect 60028 -83828 60038 -82682
rect 60092 -83828 60102 -82682
rect 60202 -83828 60212 -82682
rect 60266 -83828 60276 -82682
rect 60380 -83832 60390 -82686
rect 60444 -83832 60454 -82686
rect 60562 -83832 60572 -82686
rect 60626 -83832 60636 -82686
rect 60742 -83824 60752 -82678
rect 60806 -83824 60816 -82678
rect 60918 -83828 60928 -82682
rect 60982 -83828 60992 -82682
rect 61096 -83828 61106 -82682
rect 61160 -83828 61170 -82682
rect 61272 -83832 61282 -82686
rect 61336 -83832 61346 -82686
rect 61452 -83826 61462 -82680
rect 61516 -83826 61526 -82680
rect 61630 -83824 61640 -82678
rect 61694 -83824 61704 -82678
rect 61802 -83828 61812 -82682
rect 61866 -83828 61876 -82682
rect 61982 -83828 61992 -82682
rect 62046 -83828 62056 -82682
rect 62162 -83828 62172 -82682
rect 62226 -83828 62236 -82682
rect 62342 -83828 62352 -82682
rect 62406 -83828 62416 -82682
rect 62520 -83826 62530 -82680
rect 62584 -83826 62594 -82680
rect 62694 -83822 62704 -82676
rect 62758 -83822 62768 -82676
rect 62872 -83828 62882 -82682
rect 62936 -83828 62946 -82682
rect 63054 -83826 63064 -82680
rect 63118 -83826 63128 -82680
rect 63230 -83822 63240 -82676
rect 63294 -83822 63304 -82676
rect 63406 -83826 63416 -82680
rect 63470 -83826 63480 -82680
rect 63586 -83824 63596 -82678
rect 63650 -83824 63660 -82678
rect 63764 -83824 63774 -82678
rect 63828 -83824 63838 -82678
rect 63942 -83822 63952 -82676
rect 64006 -83822 64016 -82676
rect 64120 -83820 64130 -82674
rect 64184 -83820 64194 -82674
rect 64296 -83824 64306 -82678
rect 64360 -83824 64370 -82678
rect 56018 -84564 56312 -84342
rect 56276 -86180 56286 -85034
rect 56340 -86180 56350 -85034
rect 56452 -86178 56462 -85032
rect 56516 -86178 56526 -85032
rect 56630 -86182 56640 -85036
rect 56694 -86182 56704 -85036
rect 56814 -86178 56824 -85032
rect 56878 -86178 56888 -85032
rect 56988 -86186 56998 -85040
rect 57052 -86186 57062 -85040
rect 57164 -86190 57174 -85044
rect 57228 -86190 57238 -85044
rect 57344 -86186 57354 -85040
rect 57408 -86186 57418 -85040
rect 57520 -86182 57530 -85036
rect 57584 -86182 57594 -85036
rect 57702 -86182 57712 -85036
rect 57766 -86182 57776 -85036
rect 57878 -86186 57888 -85040
rect 57942 -86186 57952 -85040
rect 58056 -86186 58066 -85040
rect 58120 -86186 58130 -85040
rect 58238 -86190 58248 -85044
rect 58302 -86190 58312 -85044
rect 58412 -86186 58422 -85040
rect 58476 -86186 58486 -85040
rect 58592 -86184 58602 -85038
rect 58656 -86184 58666 -85038
rect 58768 -86184 58778 -85038
rect 58832 -86184 58842 -85038
rect 58948 -86182 58958 -85036
rect 59012 -86182 59022 -85036
rect 59128 -86182 59138 -85036
rect 59192 -86182 59202 -85036
rect 59306 -86182 59316 -85036
rect 59370 -86182 59380 -85036
rect 59484 -86178 59494 -85032
rect 59548 -86178 59558 -85032
rect 59660 -86182 59670 -85036
rect 59724 -86182 59734 -85036
rect 59838 -86186 59848 -85040
rect 59902 -86186 59912 -85040
rect 60016 -86186 60026 -85040
rect 60080 -86186 60090 -85040
rect 60190 -86186 60200 -85040
rect 60254 -86186 60264 -85040
rect 60368 -86190 60378 -85044
rect 60432 -86190 60442 -85044
rect 60550 -86190 60560 -85044
rect 60614 -86190 60624 -85044
rect 60730 -86182 60740 -85036
rect 60794 -86182 60804 -85036
rect 60906 -86186 60916 -85040
rect 60970 -86186 60980 -85040
rect 61084 -86186 61094 -85040
rect 61148 -86186 61158 -85040
rect 61260 -86190 61270 -85044
rect 61324 -86190 61334 -85044
rect 61440 -86184 61450 -85038
rect 61504 -86184 61514 -85038
rect 61618 -86182 61628 -85036
rect 61682 -86182 61692 -85036
rect 61790 -86186 61800 -85040
rect 61854 -86186 61864 -85040
rect 61970 -86186 61980 -85040
rect 62034 -86186 62044 -85040
rect 62150 -86186 62160 -85040
rect 62214 -86186 62224 -85040
rect 62330 -86186 62340 -85040
rect 62394 -86186 62404 -85040
rect 62508 -86184 62518 -85038
rect 62572 -86184 62582 -85038
rect 62682 -86180 62692 -85034
rect 62746 -86180 62756 -85034
rect 62860 -86186 62870 -85040
rect 62924 -86186 62934 -85040
rect 63042 -86184 63052 -85038
rect 63106 -86184 63116 -85038
rect 63218 -86180 63228 -85034
rect 63282 -86180 63292 -85034
rect 63394 -86184 63404 -85038
rect 63458 -86184 63468 -85038
rect 63574 -86182 63584 -85036
rect 63638 -86182 63648 -85036
rect 63752 -86182 63762 -85036
rect 63816 -86182 63826 -85036
rect 63930 -86180 63940 -85034
rect 63994 -86180 64004 -85034
rect 64108 -86178 64118 -85032
rect 64172 -86178 64182 -85032
rect 64284 -86182 64294 -85036
rect 64348 -86182 64358 -85036
rect 56326 -86428 56336 -86272
rect 56442 -86428 56452 -86272
rect 56508 -86434 56518 -86278
rect 56624 -86434 56634 -86278
rect 56690 -86430 56700 -86274
rect 56806 -86430 56816 -86274
rect 56870 -86430 56880 -86274
rect 56986 -86430 56996 -86274
rect 57048 -86428 57058 -86272
rect 57164 -86428 57174 -86272
rect 57224 -86428 57234 -86272
rect 57340 -86428 57350 -86272
rect 57408 -86430 57418 -86274
rect 57524 -86430 57534 -86274
rect 57582 -86430 57592 -86274
rect 57698 -86430 57708 -86274
rect 57756 -86430 57766 -86274
rect 57872 -86430 57882 -86274
rect 57938 -86434 57948 -86278
rect 58054 -86434 58064 -86278
rect 58112 -86430 58122 -86274
rect 58228 -86430 58238 -86274
rect 58290 -86430 58300 -86274
rect 58406 -86430 58416 -86274
rect 58470 -86430 58480 -86274
rect 58586 -86430 58596 -86274
rect 58640 -86430 58650 -86274
rect 58756 -86430 58766 -86274
rect 58820 -86430 58830 -86274
rect 58936 -86430 58946 -86274
rect 59004 -86430 59014 -86274
rect 59120 -86430 59130 -86274
rect 59178 -86430 59188 -86274
rect 59294 -86430 59304 -86274
rect 59352 -86428 59362 -86272
rect 59468 -86428 59478 -86272
rect 59530 -86424 59540 -86268
rect 59646 -86424 59656 -86268
rect 59712 -86434 59722 -86278
rect 59828 -86434 59838 -86278
rect 59888 -86430 59898 -86274
rect 60004 -86430 60014 -86274
rect 60068 -86430 60078 -86274
rect 60184 -86430 60194 -86274
rect 60240 -86430 60250 -86274
rect 60356 -86430 60366 -86274
rect 60424 -86434 60434 -86278
rect 60540 -86434 60550 -86278
rect 60598 -86430 60608 -86274
rect 60714 -86430 60724 -86274
rect 60778 -86434 60788 -86278
rect 60894 -86434 60904 -86278
rect 60954 -86434 60964 -86278
rect 61070 -86434 61080 -86278
rect 61130 -86430 61140 -86274
rect 61246 -86430 61256 -86274
rect 61310 -86434 61320 -86278
rect 61426 -86434 61436 -86278
rect 61490 -86430 61500 -86274
rect 61606 -86430 61616 -86274
rect 61668 -86438 61678 -86282
rect 61784 -86438 61794 -86282
rect 61848 -86430 61858 -86274
rect 61964 -86430 61974 -86274
rect 62024 -86434 62034 -86278
rect 62140 -86434 62150 -86278
rect 62202 -86424 62212 -86268
rect 62318 -86424 62328 -86268
rect 62380 -86430 62390 -86274
rect 62496 -86430 62506 -86274
rect 62558 -86430 62568 -86274
rect 62674 -86430 62684 -86274
rect 62738 -86434 62748 -86278
rect 62854 -86434 62864 -86278
rect 62918 -86434 62928 -86278
rect 63034 -86434 63044 -86278
rect 63092 -86430 63102 -86274
rect 63208 -86430 63218 -86274
rect 63276 -86434 63286 -86278
rect 63392 -86434 63402 -86278
rect 63444 -86434 63454 -86278
rect 63560 -86434 63570 -86278
rect 63622 -86440 63632 -86284
rect 63738 -86440 63748 -86284
rect 63810 -86428 63820 -86272
rect 63926 -86428 63936 -86272
rect 63982 -86430 63992 -86274
rect 64098 -86430 64108 -86274
rect 64162 -86428 64172 -86272
rect 64278 -86428 64288 -86272
rect 56260 -87642 56270 -86496
rect 56324 -87642 56334 -86496
rect 56436 -87640 56446 -86494
rect 56500 -87640 56510 -86494
rect 56614 -87644 56624 -86498
rect 56678 -87644 56688 -86498
rect 56798 -87640 56808 -86494
rect 56862 -87640 56872 -86494
rect 56972 -87648 56982 -86502
rect 57036 -87648 57046 -86502
rect 57148 -87652 57158 -86506
rect 57212 -87652 57222 -86506
rect 57328 -87648 57338 -86502
rect 57392 -87648 57402 -86502
rect 57504 -87644 57514 -86498
rect 57568 -87644 57578 -86498
rect 57686 -87644 57696 -86498
rect 57750 -87644 57760 -86498
rect 57862 -87648 57872 -86502
rect 57926 -87648 57936 -86502
rect 58040 -87648 58050 -86502
rect 58104 -87648 58114 -86502
rect 58222 -87652 58232 -86506
rect 58286 -87652 58296 -86506
rect 58396 -87648 58406 -86502
rect 58460 -87648 58470 -86502
rect 58576 -87646 58586 -86500
rect 58640 -87646 58650 -86500
rect 58752 -87646 58762 -86500
rect 58816 -87646 58826 -86500
rect 58932 -87644 58942 -86498
rect 58996 -87644 59006 -86498
rect 59112 -87644 59122 -86498
rect 59176 -87644 59186 -86498
rect 59290 -87644 59300 -86498
rect 59354 -87644 59364 -86498
rect 59468 -87640 59478 -86494
rect 59532 -87640 59542 -86494
rect 59644 -87644 59654 -86498
rect 59708 -87644 59718 -86498
rect 59822 -87648 59832 -86502
rect 59886 -87648 59896 -86502
rect 60000 -87648 60010 -86502
rect 60064 -87648 60074 -86502
rect 60174 -87648 60184 -86502
rect 60238 -87648 60248 -86502
rect 60352 -87652 60362 -86506
rect 60416 -87652 60426 -86506
rect 60534 -87652 60544 -86506
rect 60598 -87652 60608 -86506
rect 60714 -87644 60724 -86498
rect 60778 -87644 60788 -86498
rect 60890 -87648 60900 -86502
rect 60954 -87648 60964 -86502
rect 61068 -87648 61078 -86502
rect 61132 -87648 61142 -86502
rect 61244 -87652 61254 -86506
rect 61308 -87652 61318 -86506
rect 61424 -87646 61434 -86500
rect 61488 -87646 61498 -86500
rect 61602 -87644 61612 -86498
rect 61666 -87644 61676 -86498
rect 61774 -87648 61784 -86502
rect 61838 -87648 61848 -86502
rect 61954 -87648 61964 -86502
rect 62018 -87648 62028 -86502
rect 62134 -87648 62144 -86502
rect 62198 -87648 62208 -86502
rect 62314 -87648 62324 -86502
rect 62378 -87648 62388 -86502
rect 62492 -87646 62502 -86500
rect 62556 -87646 62566 -86500
rect 62666 -87642 62676 -86496
rect 62730 -87642 62740 -86496
rect 62844 -87648 62854 -86502
rect 62908 -87648 62918 -86502
rect 63026 -87646 63036 -86500
rect 63090 -87646 63100 -86500
rect 63202 -87642 63212 -86496
rect 63266 -87642 63276 -86496
rect 63378 -87646 63388 -86500
rect 63442 -87646 63452 -86500
rect 63558 -87644 63568 -86498
rect 63622 -87644 63632 -86498
rect 63736 -87644 63746 -86498
rect 63800 -87644 63810 -86498
rect 63914 -87642 63924 -86496
rect 63978 -87642 63988 -86496
rect 64092 -87640 64102 -86494
rect 64156 -87640 64166 -86494
rect 64268 -87644 64278 -86498
rect 64332 -87644 64342 -86498
rect 66130 -87790 66140 -87616
rect 66196 -87790 66206 -87616
rect 66308 -87788 66318 -87614
rect 66374 -87788 66384 -87614
rect 66488 -87786 66498 -87612
rect 66554 -87786 66564 -87612
rect 66666 -87788 66676 -87614
rect 66732 -87788 66742 -87614
rect 66838 -87788 66848 -87614
rect 66904 -87788 66914 -87614
rect 67020 -87786 67030 -87612
rect 67086 -87786 67096 -87612
rect 67198 -87786 67208 -87612
rect 67264 -87786 67274 -87612
rect 55732 -88354 55742 -87954
rect 56040 -88038 56050 -87954
rect 66202 -87990 66212 -87838
rect 66316 -87990 66326 -87838
rect 66382 -87990 66392 -87838
rect 66496 -87990 66506 -87838
rect 66560 -87990 66570 -87838
rect 66674 -87990 66684 -87838
rect 66736 -87990 66746 -87838
rect 66850 -87990 66860 -87838
rect 66914 -87990 66924 -87838
rect 67028 -87990 67038 -87838
rect 67090 -87990 67100 -87838
rect 67204 -87990 67214 -87838
rect 56040 -88060 64432 -88038
rect 56040 -88094 56400 -88060
rect 56434 -88094 56472 -88060
rect 56506 -88094 56544 -88060
rect 56578 -88094 56616 -88060
rect 56650 -88094 56688 -88060
rect 56722 -88094 56760 -88060
rect 56794 -88094 56832 -88060
rect 56866 -88094 56904 -88060
rect 56938 -88094 56976 -88060
rect 57010 -88094 57048 -88060
rect 57082 -88094 57120 -88060
rect 57154 -88094 57192 -88060
rect 57226 -88094 57264 -88060
rect 57298 -88094 57336 -88060
rect 57370 -88094 57408 -88060
rect 57442 -88094 57480 -88060
rect 57514 -88094 57552 -88060
rect 57586 -88094 57624 -88060
rect 57658 -88094 57696 -88060
rect 57730 -88094 57768 -88060
rect 57802 -88094 57840 -88060
rect 57874 -88094 57912 -88060
rect 57946 -88094 57984 -88060
rect 58018 -88094 58056 -88060
rect 58090 -88094 58128 -88060
rect 58162 -88094 58200 -88060
rect 58234 -88094 58272 -88060
rect 58306 -88094 58344 -88060
rect 58378 -88094 58416 -88060
rect 58450 -88094 58488 -88060
rect 58522 -88094 58560 -88060
rect 58594 -88094 58632 -88060
rect 58666 -88094 58704 -88060
rect 58738 -88094 58776 -88060
rect 58810 -88094 58848 -88060
rect 58882 -88094 58920 -88060
rect 58954 -88094 58992 -88060
rect 59026 -88094 59064 -88060
rect 59098 -88094 59136 -88060
rect 59170 -88094 59208 -88060
rect 59242 -88094 59280 -88060
rect 59314 -88094 59352 -88060
rect 59386 -88094 59424 -88060
rect 59458 -88094 59496 -88060
rect 59530 -88094 59568 -88060
rect 59602 -88094 59640 -88060
rect 59674 -88094 59712 -88060
rect 59746 -88094 59784 -88060
rect 59818 -88094 59856 -88060
rect 59890 -88094 59928 -88060
rect 59962 -88094 60000 -88060
rect 60034 -88094 60072 -88060
rect 60106 -88094 60144 -88060
rect 60178 -88094 60216 -88060
rect 60250 -88094 60288 -88060
rect 60322 -88094 60360 -88060
rect 60394 -88094 60432 -88060
rect 60466 -88094 60504 -88060
rect 60538 -88094 60576 -88060
rect 60610 -88094 60648 -88060
rect 60682 -88094 60720 -88060
rect 60754 -88094 60792 -88060
rect 60826 -88094 60864 -88060
rect 60898 -88094 60936 -88060
rect 60970 -88094 61008 -88060
rect 61042 -88094 61080 -88060
rect 61114 -88094 61152 -88060
rect 61186 -88094 61224 -88060
rect 61258 -88094 61296 -88060
rect 61330 -88094 61368 -88060
rect 61402 -88094 61440 -88060
rect 61474 -88094 61512 -88060
rect 61546 -88094 61584 -88060
rect 61618 -88094 61656 -88060
rect 61690 -88094 61728 -88060
rect 61762 -88094 61800 -88060
rect 61834 -88094 61872 -88060
rect 61906 -88094 61944 -88060
rect 61978 -88094 62016 -88060
rect 62050 -88094 62088 -88060
rect 62122 -88094 62160 -88060
rect 62194 -88094 62232 -88060
rect 62266 -88094 62304 -88060
rect 62338 -88094 62376 -88060
rect 62410 -88094 62448 -88060
rect 62482 -88094 62520 -88060
rect 62554 -88094 62592 -88060
rect 62626 -88094 62664 -88060
rect 62698 -88094 62736 -88060
rect 62770 -88094 62808 -88060
rect 62842 -88094 62880 -88060
rect 62914 -88094 62952 -88060
rect 62986 -88094 63024 -88060
rect 63058 -88094 63096 -88060
rect 63130 -88094 63168 -88060
rect 63202 -88094 63240 -88060
rect 63274 -88094 63312 -88060
rect 63346 -88094 63384 -88060
rect 63418 -88094 63456 -88060
rect 63490 -88094 63528 -88060
rect 63562 -88094 63600 -88060
rect 63634 -88094 63672 -88060
rect 63706 -88094 63744 -88060
rect 63778 -88094 63816 -88060
rect 63850 -88094 63888 -88060
rect 63922 -88094 63960 -88060
rect 63994 -88094 64032 -88060
rect 64066 -88094 64104 -88060
rect 64138 -88094 64176 -88060
rect 64210 -88094 64248 -88060
rect 64282 -88094 64432 -88060
rect 56040 -88134 64432 -88094
rect 56040 -88168 56400 -88134
rect 56434 -88168 56472 -88134
rect 56506 -88168 56544 -88134
rect 56578 -88168 56616 -88134
rect 56650 -88168 56688 -88134
rect 56722 -88168 56760 -88134
rect 56794 -88168 56832 -88134
rect 56866 -88168 56904 -88134
rect 56938 -88168 56976 -88134
rect 57010 -88168 57048 -88134
rect 57082 -88168 57120 -88134
rect 57154 -88168 57192 -88134
rect 57226 -88168 57264 -88134
rect 57298 -88168 57336 -88134
rect 57370 -88168 57408 -88134
rect 57442 -88168 57480 -88134
rect 57514 -88168 57552 -88134
rect 57586 -88168 57624 -88134
rect 57658 -88168 57696 -88134
rect 57730 -88168 57768 -88134
rect 57802 -88168 57840 -88134
rect 57874 -88168 57912 -88134
rect 57946 -88168 57984 -88134
rect 58018 -88168 58056 -88134
rect 58090 -88168 58128 -88134
rect 58162 -88168 58200 -88134
rect 58234 -88168 58272 -88134
rect 58306 -88168 58344 -88134
rect 58378 -88168 58416 -88134
rect 58450 -88168 58488 -88134
rect 58522 -88168 58560 -88134
rect 58594 -88168 58632 -88134
rect 58666 -88168 58704 -88134
rect 58738 -88168 58776 -88134
rect 58810 -88168 58848 -88134
rect 58882 -88168 58920 -88134
rect 58954 -88168 58992 -88134
rect 59026 -88168 59064 -88134
rect 59098 -88168 59136 -88134
rect 59170 -88168 59208 -88134
rect 59242 -88168 59280 -88134
rect 59314 -88168 59352 -88134
rect 59386 -88168 59424 -88134
rect 59458 -88168 59496 -88134
rect 59530 -88168 59568 -88134
rect 59602 -88168 59640 -88134
rect 59674 -88168 59712 -88134
rect 59746 -88168 59784 -88134
rect 59818 -88168 59856 -88134
rect 59890 -88168 59928 -88134
rect 59962 -88168 60000 -88134
rect 60034 -88168 60072 -88134
rect 60106 -88168 60144 -88134
rect 60178 -88168 60216 -88134
rect 60250 -88168 60288 -88134
rect 60322 -88168 60360 -88134
rect 60394 -88168 60432 -88134
rect 60466 -88168 60504 -88134
rect 60538 -88168 60576 -88134
rect 60610 -88168 60648 -88134
rect 60682 -88168 60720 -88134
rect 60754 -88168 60792 -88134
rect 60826 -88168 60864 -88134
rect 60898 -88168 60936 -88134
rect 60970 -88168 61008 -88134
rect 61042 -88168 61080 -88134
rect 61114 -88168 61152 -88134
rect 61186 -88168 61224 -88134
rect 61258 -88168 61296 -88134
rect 61330 -88168 61368 -88134
rect 61402 -88168 61440 -88134
rect 61474 -88168 61512 -88134
rect 61546 -88168 61584 -88134
rect 61618 -88168 61656 -88134
rect 61690 -88168 61728 -88134
rect 61762 -88168 61800 -88134
rect 61834 -88168 61872 -88134
rect 61906 -88168 61944 -88134
rect 61978 -88168 62016 -88134
rect 62050 -88168 62088 -88134
rect 62122 -88168 62160 -88134
rect 62194 -88168 62232 -88134
rect 62266 -88168 62304 -88134
rect 62338 -88168 62376 -88134
rect 62410 -88168 62448 -88134
rect 62482 -88168 62520 -88134
rect 62554 -88168 62592 -88134
rect 62626 -88168 62664 -88134
rect 62698 -88168 62736 -88134
rect 62770 -88168 62808 -88134
rect 62842 -88168 62880 -88134
rect 62914 -88168 62952 -88134
rect 62986 -88168 63024 -88134
rect 63058 -88168 63096 -88134
rect 63130 -88168 63168 -88134
rect 63202 -88168 63240 -88134
rect 63274 -88168 63312 -88134
rect 63346 -88168 63384 -88134
rect 63418 -88168 63456 -88134
rect 63490 -88168 63528 -88134
rect 63562 -88168 63600 -88134
rect 63634 -88168 63672 -88134
rect 63706 -88168 63744 -88134
rect 63778 -88168 63816 -88134
rect 63850 -88168 63888 -88134
rect 63922 -88168 63960 -88134
rect 63994 -88168 64032 -88134
rect 64066 -88168 64104 -88134
rect 64138 -88168 64176 -88134
rect 64210 -88168 64248 -88134
rect 64282 -88168 64432 -88134
rect 56040 -88208 64432 -88168
rect 56040 -88242 56400 -88208
rect 56434 -88242 56472 -88208
rect 56506 -88242 56544 -88208
rect 56578 -88242 56616 -88208
rect 56650 -88242 56688 -88208
rect 56722 -88242 56760 -88208
rect 56794 -88242 56832 -88208
rect 56866 -88242 56904 -88208
rect 56938 -88242 56976 -88208
rect 57010 -88242 57048 -88208
rect 57082 -88242 57120 -88208
rect 57154 -88242 57192 -88208
rect 57226 -88242 57264 -88208
rect 57298 -88242 57336 -88208
rect 57370 -88242 57408 -88208
rect 57442 -88242 57480 -88208
rect 57514 -88242 57552 -88208
rect 57586 -88242 57624 -88208
rect 57658 -88242 57696 -88208
rect 57730 -88242 57768 -88208
rect 57802 -88242 57840 -88208
rect 57874 -88242 57912 -88208
rect 57946 -88242 57984 -88208
rect 58018 -88242 58056 -88208
rect 58090 -88242 58128 -88208
rect 58162 -88242 58200 -88208
rect 58234 -88242 58272 -88208
rect 58306 -88242 58344 -88208
rect 58378 -88242 58416 -88208
rect 58450 -88242 58488 -88208
rect 58522 -88242 58560 -88208
rect 58594 -88242 58632 -88208
rect 58666 -88242 58704 -88208
rect 58738 -88242 58776 -88208
rect 58810 -88242 58848 -88208
rect 58882 -88242 58920 -88208
rect 58954 -88242 58992 -88208
rect 59026 -88242 59064 -88208
rect 59098 -88242 59136 -88208
rect 59170 -88242 59208 -88208
rect 59242 -88242 59280 -88208
rect 59314 -88242 59352 -88208
rect 59386 -88242 59424 -88208
rect 59458 -88242 59496 -88208
rect 59530 -88242 59568 -88208
rect 59602 -88242 59640 -88208
rect 59674 -88242 59712 -88208
rect 59746 -88242 59784 -88208
rect 59818 -88242 59856 -88208
rect 59890 -88242 59928 -88208
rect 59962 -88242 60000 -88208
rect 60034 -88242 60072 -88208
rect 60106 -88242 60144 -88208
rect 60178 -88242 60216 -88208
rect 60250 -88242 60288 -88208
rect 60322 -88242 60360 -88208
rect 60394 -88242 60432 -88208
rect 60466 -88242 60504 -88208
rect 60538 -88242 60576 -88208
rect 60610 -88242 60648 -88208
rect 60682 -88242 60720 -88208
rect 60754 -88242 60792 -88208
rect 60826 -88242 60864 -88208
rect 60898 -88242 60936 -88208
rect 60970 -88242 61008 -88208
rect 61042 -88242 61080 -88208
rect 61114 -88242 61152 -88208
rect 61186 -88242 61224 -88208
rect 61258 -88242 61296 -88208
rect 61330 -88242 61368 -88208
rect 61402 -88242 61440 -88208
rect 61474 -88242 61512 -88208
rect 61546 -88242 61584 -88208
rect 61618 -88242 61656 -88208
rect 61690 -88242 61728 -88208
rect 61762 -88242 61800 -88208
rect 61834 -88242 61872 -88208
rect 61906 -88242 61944 -88208
rect 61978 -88242 62016 -88208
rect 62050 -88242 62088 -88208
rect 62122 -88242 62160 -88208
rect 62194 -88242 62232 -88208
rect 62266 -88242 62304 -88208
rect 62338 -88242 62376 -88208
rect 62410 -88242 62448 -88208
rect 62482 -88242 62520 -88208
rect 62554 -88242 62592 -88208
rect 62626 -88242 62664 -88208
rect 62698 -88242 62736 -88208
rect 62770 -88242 62808 -88208
rect 62842 -88242 62880 -88208
rect 62914 -88242 62952 -88208
rect 62986 -88242 63024 -88208
rect 63058 -88242 63096 -88208
rect 63130 -88242 63168 -88208
rect 63202 -88242 63240 -88208
rect 63274 -88242 63312 -88208
rect 63346 -88242 63384 -88208
rect 63418 -88242 63456 -88208
rect 63490 -88242 63528 -88208
rect 63562 -88242 63600 -88208
rect 63634 -88242 63672 -88208
rect 63706 -88242 63744 -88208
rect 63778 -88242 63816 -88208
rect 63850 -88242 63888 -88208
rect 63922 -88242 63960 -88208
rect 63994 -88242 64032 -88208
rect 64066 -88242 64104 -88208
rect 64138 -88242 64176 -88208
rect 64210 -88242 64248 -88208
rect 64282 -88242 64432 -88208
rect 66136 -88218 66146 -88044
rect 66202 -88218 66212 -88044
rect 66316 -88214 66326 -88040
rect 66382 -88214 66392 -88040
rect 66496 -88216 66506 -88042
rect 66562 -88216 66572 -88042
rect 66674 -88216 66684 -88042
rect 66740 -88216 66750 -88042
rect 66852 -88216 66862 -88042
rect 66918 -88216 66928 -88042
rect 67030 -88216 67040 -88042
rect 67096 -88216 67106 -88042
rect 67208 -88220 67218 -88046
rect 67274 -88220 67284 -88046
rect 56040 -88292 64432 -88242
rect 56040 -88354 56050 -88292
rect 54844 -89048 65498 -88612
rect 66126 -88626 66136 -88452
rect 66192 -88626 66202 -88452
rect 66310 -88620 66320 -88446
rect 66376 -88620 66386 -88446
rect 66490 -88624 66500 -88450
rect 66556 -88624 66566 -88450
rect 66666 -88626 66676 -88452
rect 66732 -88626 66742 -88452
rect 66844 -88620 66854 -88446
rect 66910 -88620 66920 -88446
rect 67024 -88622 67034 -88448
rect 67090 -88622 67100 -88448
rect 67202 -88626 67212 -88452
rect 67268 -88626 67278 -88452
rect 66200 -88826 66210 -88674
rect 66314 -88826 66324 -88674
rect 66382 -88828 66392 -88676
rect 66496 -88828 66506 -88676
rect 66554 -88830 66564 -88678
rect 66668 -88830 66678 -88678
rect 66736 -88830 66746 -88678
rect 66850 -88830 66860 -88678
rect 66914 -88830 66924 -88678
rect 67028 -88830 67038 -88678
rect 67094 -88830 67104 -88678
rect 67208 -88830 67218 -88678
rect 66130 -89028 66140 -88874
rect 66192 -89028 66202 -88874
rect 66310 -89034 66320 -88880
rect 66372 -89034 66382 -88880
rect 66486 -89030 66496 -88876
rect 66548 -89030 66558 -88876
rect 66662 -89034 66672 -88880
rect 66724 -89034 66734 -88880
rect 66842 -89036 66852 -88882
rect 66904 -89036 66914 -88882
rect 67024 -89034 67034 -88880
rect 67086 -89034 67096 -88880
rect 67214 -89036 67224 -88882
rect 67276 -89036 67286 -88882
rect 68250 -89018 68260 -87882
rect 68312 -89018 68322 -87882
rect 68432 -89012 68442 -87876
rect 68494 -89012 68504 -87876
rect 68618 -89020 68628 -87884
rect 68680 -89020 68690 -87884
rect 68792 -89026 68802 -87890
rect 68854 -89026 68864 -87890
rect 68970 -89026 68980 -87890
rect 69032 -89026 69042 -87890
rect 69150 -89026 69160 -87890
rect 69212 -89026 69222 -87890
rect 69326 -89026 69336 -87890
rect 69388 -89026 69398 -87890
rect 69504 -89022 69514 -87886
rect 69566 -89022 69576 -87886
rect 69684 -89024 69694 -87888
rect 69746 -89024 69756 -87888
rect 69858 -89022 69868 -87886
rect 69920 -89022 69930 -87886
rect 70038 -89026 70048 -87890
rect 70100 -89026 70110 -87890
rect 70214 -89024 70224 -87888
rect 70276 -89024 70286 -87888
rect 70394 -89024 70404 -87888
rect 70456 -89024 70466 -87888
rect 70572 -89026 70582 -87890
rect 70634 -89026 70644 -87890
rect 70750 -89028 70760 -87892
rect 70812 -89028 70822 -87892
rect 70926 -89026 70936 -87890
rect 70988 -89026 70998 -87890
rect 71104 -89028 71114 -87892
rect 71166 -89028 71176 -87892
rect 71284 -89026 71294 -87890
rect 71346 -89026 71356 -87890
rect 71462 -89026 71472 -87890
rect 71524 -89026 71534 -87890
rect 71638 -89028 71648 -87892
rect 71700 -89028 71710 -87892
rect 71816 -89026 71826 -87890
rect 71878 -89026 71888 -87890
rect 56408 -89246 56418 -89192
rect 56534 -89246 56544 -89192
rect 56588 -89248 56598 -89194
rect 56714 -89248 56724 -89194
rect 56774 -89248 56784 -89194
rect 56900 -89248 56910 -89194
rect 56958 -89246 56968 -89192
rect 57084 -89246 57094 -89192
rect 57134 -89246 57144 -89192
rect 57260 -89246 57270 -89192
rect 57308 -89246 57318 -89192
rect 57434 -89246 57444 -89192
rect 57484 -89248 57494 -89194
rect 57610 -89248 57620 -89194
rect 57672 -89254 57682 -89200
rect 57798 -89254 57808 -89200
rect 57846 -89254 57856 -89200
rect 57972 -89254 57982 -89200
rect 58028 -89266 58038 -89212
rect 58154 -89266 58164 -89212
rect 58204 -89268 58214 -89210
rect 58292 -89268 58302 -89210
rect 58402 -89266 58412 -89208
rect 58490 -89266 58500 -89208
rect 58564 -89266 58574 -89208
rect 58652 -89266 58662 -89208
rect 58750 -89266 58760 -89208
rect 58838 -89266 58848 -89208
rect 58926 -89268 58936 -89210
rect 59014 -89268 59024 -89210
rect 59098 -89266 59108 -89208
rect 59186 -89266 59196 -89208
rect 59282 -89266 59292 -89208
rect 59370 -89266 59380 -89208
rect 59458 -89262 59468 -89204
rect 59546 -89262 59556 -89204
rect 59632 -89262 59642 -89204
rect 59720 -89262 59730 -89204
rect 59822 -89266 59832 -89208
rect 59910 -89266 59920 -89208
rect 60864 -89262 60874 -89204
rect 60952 -89262 60962 -89204
rect 61054 -89266 61064 -89208
rect 61142 -89266 61152 -89208
rect 61232 -89268 61242 -89210
rect 61320 -89268 61330 -89210
rect 61406 -89262 61416 -89204
rect 61494 -89262 61504 -89204
rect 61584 -89254 61594 -89196
rect 61672 -89254 61682 -89196
rect 61760 -89262 61770 -89204
rect 61848 -89262 61858 -89204
rect 61952 -89262 61962 -89204
rect 62040 -89262 62050 -89204
rect 62112 -89258 62122 -89200
rect 62200 -89258 62210 -89200
rect 62288 -89262 62298 -89204
rect 62376 -89262 62386 -89204
rect 62468 -89262 62478 -89204
rect 62556 -89262 62566 -89204
rect 62642 -89266 62652 -89208
rect 62730 -89266 62740 -89208
rect 62832 -89258 62842 -89200
rect 62920 -89258 62930 -89200
rect 63016 -89258 63026 -89200
rect 63104 -89258 63114 -89200
rect 63178 -89258 63188 -89200
rect 63266 -89258 63276 -89200
rect 63360 -89262 63370 -89204
rect 63448 -89262 63458 -89204
rect 63544 -89266 63554 -89208
rect 63632 -89266 63642 -89208
rect 63706 -89258 63716 -89200
rect 63794 -89258 63804 -89200
rect 63890 -89258 63900 -89200
rect 63978 -89258 63988 -89200
rect 64078 -89258 64088 -89200
rect 64166 -89258 64176 -89200
rect 64246 -89258 64256 -89200
rect 64334 -89258 64344 -89200
rect 56352 -90484 56362 -89326
rect 56414 -90484 56424 -89326
rect 56538 -90484 56548 -89326
rect 56600 -90484 56610 -89326
rect 56710 -90492 56720 -89334
rect 56772 -90492 56782 -89334
rect 56896 -90484 56906 -89326
rect 56958 -90484 56968 -89326
rect 57062 -90484 57072 -89326
rect 57124 -90484 57134 -89326
rect 57250 -90484 57260 -89326
rect 57312 -90484 57322 -89326
rect 57424 -90486 57434 -89328
rect 57486 -90486 57496 -89328
rect 57604 -90486 57614 -89328
rect 57666 -90486 57676 -89328
rect 57770 -90486 57780 -89328
rect 57832 -90486 57842 -89328
rect 57964 -90484 57974 -89326
rect 58026 -90484 58036 -89326
rect 58132 -90476 58142 -89318
rect 58194 -90476 58204 -89318
rect 58318 -90480 58328 -89322
rect 58380 -90480 58390 -89322
rect 58490 -90484 58500 -89326
rect 58552 -90484 58562 -89326
rect 58676 -90480 58686 -89322
rect 58738 -90480 58748 -89322
rect 58848 -90484 58858 -89326
rect 58910 -90484 58920 -89326
rect 59028 -90486 59038 -89328
rect 59090 -90486 59100 -89328
rect 59204 -90488 59214 -89330
rect 59266 -90488 59276 -89330
rect 59386 -90486 59396 -89328
rect 59448 -90486 59458 -89328
rect 59560 -90484 59570 -89326
rect 59622 -90484 59632 -89326
rect 59742 -90484 59752 -89326
rect 59804 -90484 59814 -89326
rect 59912 -90480 59922 -89322
rect 59974 -90480 59984 -89322
rect 60786 -90484 60796 -89326
rect 60848 -90484 60858 -89326
rect 60970 -90484 60980 -89326
rect 61032 -90484 61042 -89326
rect 61132 -90484 61142 -89326
rect 61194 -90484 61204 -89326
rect 61320 -90486 61330 -89328
rect 61382 -90486 61392 -89328
rect 61496 -90486 61506 -89328
rect 61558 -90486 61568 -89328
rect 61680 -90486 61690 -89328
rect 61742 -90486 61752 -89328
rect 61852 -90490 61862 -89332
rect 61914 -90490 61924 -89332
rect 62032 -90484 62042 -89326
rect 62094 -90484 62104 -89326
rect 62206 -90480 62216 -89322
rect 62268 -90480 62278 -89322
rect 62388 -90484 62398 -89326
rect 62450 -90484 62460 -89326
rect 62560 -90480 62570 -89322
rect 62622 -90480 62632 -89322
rect 62746 -90484 62756 -89326
rect 62808 -90484 62818 -89326
rect 62916 -90484 62926 -89326
rect 62978 -90484 62988 -89326
rect 63102 -90478 63112 -89320
rect 63164 -90478 63174 -89320
rect 63278 -90480 63288 -89322
rect 63340 -90480 63350 -89322
rect 63458 -90486 63468 -89328
rect 63520 -90486 63530 -89328
rect 63628 -90490 63638 -89332
rect 63690 -90490 63700 -89332
rect 63816 -90484 63826 -89326
rect 63878 -90484 63888 -89326
rect 63984 -90486 63994 -89328
rect 64046 -90486 64056 -89328
rect 64174 -90484 64184 -89326
rect 64236 -90484 64246 -89326
rect 64338 -90486 64348 -89328
rect 64400 -90486 64410 -89328
rect 64592 -89678 65456 -89048
rect 68320 -89228 68330 -89082
rect 68424 -89228 68434 -89082
rect 68500 -89228 68510 -89082
rect 68604 -89228 68614 -89082
rect 68680 -89228 68690 -89082
rect 68784 -89228 68794 -89082
rect 68858 -89228 68868 -89082
rect 68962 -89228 68972 -89082
rect 69034 -89228 69044 -89082
rect 69138 -89228 69148 -89082
rect 69214 -89230 69224 -89084
rect 69318 -89230 69328 -89084
rect 69390 -89228 69400 -89082
rect 69494 -89228 69504 -89082
rect 69568 -89228 69578 -89082
rect 69672 -89228 69682 -89082
rect 69750 -89228 69760 -89082
rect 69854 -89228 69864 -89082
rect 69924 -89226 69934 -89080
rect 70028 -89226 70038 -89080
rect 70104 -89228 70114 -89082
rect 70208 -89228 70218 -89082
rect 70280 -89230 70290 -89084
rect 70384 -89230 70394 -89084
rect 70460 -89228 70470 -89082
rect 70564 -89228 70574 -89082
rect 70634 -89226 70644 -89080
rect 70738 -89226 70748 -89080
rect 70814 -89224 70824 -89078
rect 70918 -89224 70928 -89078
rect 70992 -89228 71002 -89082
rect 71096 -89228 71106 -89082
rect 71170 -89226 71180 -89080
rect 71274 -89226 71284 -89080
rect 71350 -89228 71360 -89082
rect 71454 -89228 71464 -89082
rect 71526 -89228 71536 -89082
rect 71630 -89228 71640 -89082
rect 71704 -89228 71714 -89082
rect 71808 -89228 71818 -89082
rect 68258 -90444 68268 -89308
rect 68320 -90444 68330 -89308
rect 68436 -90444 68446 -89308
rect 68498 -90444 68508 -89308
rect 68610 -90442 68620 -89306
rect 68672 -90442 68682 -89306
rect 68792 -90446 68802 -89310
rect 68854 -90446 68864 -89310
rect 68970 -90444 68980 -89308
rect 69032 -90444 69042 -89308
rect 69146 -90442 69156 -89306
rect 69208 -90442 69218 -89306
rect 69324 -90446 69334 -89310
rect 69386 -90446 69396 -89310
rect 69502 -90444 69512 -89308
rect 69564 -90444 69574 -89308
rect 69680 -90442 69690 -89306
rect 69742 -90442 69752 -89306
rect 69856 -90446 69866 -89310
rect 69918 -90446 69928 -89310
rect 70036 -90444 70046 -89308
rect 70098 -90444 70108 -89308
rect 70216 -90444 70226 -89308
rect 70278 -90444 70288 -89308
rect 70396 -90444 70406 -89308
rect 70458 -90444 70468 -89308
rect 70570 -90444 70580 -89308
rect 70632 -90444 70642 -89308
rect 70748 -90442 70758 -89306
rect 70810 -90442 70820 -89306
rect 70924 -90442 70934 -89306
rect 70986 -90442 70996 -89306
rect 71104 -90442 71114 -89306
rect 71166 -90442 71176 -89306
rect 71282 -90448 71292 -89312
rect 71344 -90448 71354 -89312
rect 71462 -90444 71472 -89308
rect 71524 -90444 71534 -89308
rect 71638 -90446 71648 -89310
rect 71700 -90446 71710 -89310
rect 71816 -90446 71826 -89310
rect 71878 -90446 71888 -89310
rect 72130 -91190 73922 -87728
rect 74146 -89016 74156 -87880
rect 74208 -89016 74218 -87880
rect 74328 -89010 74338 -87874
rect 74390 -89010 74400 -87874
rect 74514 -89018 74524 -87882
rect 74576 -89018 74586 -87882
rect 74688 -89024 74698 -87888
rect 74750 -89024 74760 -87888
rect 74866 -89024 74876 -87888
rect 74928 -89024 74938 -87888
rect 75046 -89024 75056 -87888
rect 75108 -89024 75118 -87888
rect 75222 -89024 75232 -87888
rect 75284 -89024 75294 -87888
rect 75400 -89020 75410 -87884
rect 75462 -89020 75472 -87884
rect 75580 -89022 75590 -87886
rect 75642 -89022 75652 -87886
rect 75754 -89020 75764 -87884
rect 75816 -89020 75826 -87884
rect 75934 -89024 75944 -87888
rect 75996 -89024 76006 -87888
rect 76110 -89022 76120 -87886
rect 76172 -89022 76182 -87886
rect 76290 -89022 76300 -87886
rect 76352 -89022 76362 -87886
rect 76468 -89024 76478 -87888
rect 76530 -89024 76540 -87888
rect 76646 -89026 76656 -87890
rect 76708 -89026 76718 -87890
rect 76822 -89024 76832 -87888
rect 76884 -89024 76894 -87888
rect 77000 -89026 77010 -87890
rect 77062 -89026 77072 -87890
rect 77180 -89024 77190 -87888
rect 77242 -89024 77252 -87888
rect 77358 -89024 77368 -87888
rect 77420 -89024 77430 -87888
rect 77534 -89026 77544 -87890
rect 77596 -89026 77606 -87890
rect 77712 -89024 77722 -87888
rect 77774 -89024 77784 -87888
rect 74216 -89226 74226 -89080
rect 74320 -89226 74330 -89080
rect 74396 -89226 74406 -89080
rect 74500 -89226 74510 -89080
rect 74576 -89226 74586 -89080
rect 74680 -89226 74690 -89080
rect 74754 -89226 74764 -89080
rect 74858 -89226 74868 -89080
rect 74930 -89226 74940 -89080
rect 75034 -89226 75044 -89080
rect 75110 -89228 75120 -89082
rect 75214 -89228 75224 -89082
rect 75286 -89226 75296 -89080
rect 75390 -89226 75400 -89080
rect 75464 -89226 75474 -89080
rect 75568 -89226 75578 -89080
rect 75646 -89226 75656 -89080
rect 75750 -89226 75760 -89080
rect 75820 -89224 75830 -89078
rect 75924 -89224 75934 -89078
rect 76000 -89226 76010 -89080
rect 76104 -89226 76114 -89080
rect 76176 -89228 76186 -89082
rect 76280 -89228 76290 -89082
rect 76356 -89226 76366 -89080
rect 76460 -89226 76470 -89080
rect 76530 -89224 76540 -89078
rect 76634 -89224 76644 -89078
rect 76710 -89222 76720 -89076
rect 76814 -89222 76824 -89076
rect 76888 -89226 76898 -89080
rect 76992 -89226 77002 -89080
rect 77066 -89224 77076 -89078
rect 77170 -89224 77180 -89078
rect 77246 -89226 77256 -89080
rect 77350 -89226 77360 -89080
rect 77422 -89226 77432 -89080
rect 77526 -89226 77536 -89080
rect 77600 -89226 77610 -89080
rect 77704 -89226 77714 -89080
rect 74154 -90442 74164 -89306
rect 74216 -90442 74226 -89306
rect 74332 -90442 74342 -89306
rect 74394 -90442 74404 -89306
rect 74506 -90440 74516 -89304
rect 74568 -90440 74578 -89304
rect 74688 -90444 74698 -89308
rect 74750 -90444 74760 -89308
rect 74866 -90442 74876 -89306
rect 74928 -90442 74938 -89306
rect 75042 -90440 75052 -89304
rect 75104 -90440 75114 -89304
rect 75220 -90444 75230 -89308
rect 75282 -90444 75292 -89308
rect 75398 -90442 75408 -89306
rect 75460 -90442 75470 -89306
rect 75576 -90440 75586 -89304
rect 75638 -90440 75648 -89304
rect 75752 -90444 75762 -89308
rect 75814 -90444 75824 -89308
rect 75932 -90442 75942 -89306
rect 75994 -90442 76004 -89306
rect 76112 -90442 76122 -89306
rect 76174 -90442 76184 -89306
rect 76292 -90442 76302 -89306
rect 76354 -90442 76364 -89306
rect 76466 -90442 76476 -89306
rect 76528 -90442 76538 -89306
rect 76644 -90440 76654 -89304
rect 76706 -90440 76716 -89304
rect 76820 -90440 76830 -89304
rect 76882 -90440 76892 -89304
rect 77000 -90440 77010 -89304
rect 77062 -90440 77072 -89304
rect 77178 -90446 77188 -89310
rect 77240 -90446 77250 -89310
rect 77358 -90442 77368 -89306
rect 77420 -90442 77430 -89306
rect 77534 -90444 77544 -89308
rect 77596 -90444 77606 -89308
rect 77712 -90444 77722 -89308
rect 77774 -90444 77784 -89308
rect 78098 -91190 79890 -87714
rect 80260 -89010 80270 -87874
rect 80322 -89010 80332 -87874
rect 80442 -89004 80452 -87868
rect 80504 -89004 80514 -87868
rect 80628 -89012 80638 -87876
rect 80690 -89012 80700 -87876
rect 80802 -89018 80812 -87882
rect 80864 -89018 80874 -87882
rect 80980 -89018 80990 -87882
rect 81042 -89018 81052 -87882
rect 81160 -89018 81170 -87882
rect 81222 -89018 81232 -87882
rect 81336 -89018 81346 -87882
rect 81398 -89018 81408 -87882
rect 81514 -89014 81524 -87878
rect 81576 -89014 81586 -87878
rect 81694 -89016 81704 -87880
rect 81756 -89016 81766 -87880
rect 81868 -89014 81878 -87878
rect 81930 -89014 81940 -87878
rect 82048 -89018 82058 -87882
rect 82110 -89018 82120 -87882
rect 82224 -89016 82234 -87880
rect 82286 -89016 82296 -87880
rect 82404 -89016 82414 -87880
rect 82466 -89016 82476 -87880
rect 82582 -89018 82592 -87882
rect 82644 -89018 82654 -87882
rect 82760 -89020 82770 -87884
rect 82822 -89020 82832 -87884
rect 82936 -89018 82946 -87882
rect 82998 -89018 83008 -87882
rect 83114 -89020 83124 -87884
rect 83176 -89020 83186 -87884
rect 83294 -89018 83304 -87882
rect 83356 -89018 83366 -87882
rect 83472 -89018 83482 -87882
rect 83534 -89018 83544 -87882
rect 83648 -89020 83658 -87884
rect 83710 -89020 83720 -87884
rect 83826 -89018 83836 -87882
rect 83888 -89018 83898 -87882
rect 80330 -89220 80340 -89074
rect 80434 -89220 80444 -89074
rect 80510 -89220 80520 -89074
rect 80614 -89220 80624 -89074
rect 80690 -89220 80700 -89074
rect 80794 -89220 80804 -89074
rect 80868 -89220 80878 -89074
rect 80972 -89220 80982 -89074
rect 81044 -89220 81054 -89074
rect 81148 -89220 81158 -89074
rect 81224 -89222 81234 -89076
rect 81328 -89222 81338 -89076
rect 81400 -89220 81410 -89074
rect 81504 -89220 81514 -89074
rect 81578 -89220 81588 -89074
rect 81682 -89220 81692 -89074
rect 81760 -89220 81770 -89074
rect 81864 -89220 81874 -89074
rect 81934 -89218 81944 -89072
rect 82038 -89218 82048 -89072
rect 82114 -89220 82124 -89074
rect 82218 -89220 82228 -89074
rect 82290 -89222 82300 -89076
rect 82394 -89222 82404 -89076
rect 82470 -89220 82480 -89074
rect 82574 -89220 82584 -89074
rect 82644 -89218 82654 -89072
rect 82748 -89218 82758 -89072
rect 82824 -89216 82834 -89070
rect 82928 -89216 82938 -89070
rect 83002 -89220 83012 -89074
rect 83106 -89220 83116 -89074
rect 83180 -89218 83190 -89072
rect 83284 -89218 83294 -89072
rect 83360 -89220 83370 -89074
rect 83464 -89220 83474 -89074
rect 83536 -89220 83546 -89074
rect 83640 -89220 83650 -89074
rect 83714 -89220 83724 -89074
rect 83818 -89220 83828 -89074
rect 80268 -90436 80278 -89300
rect 80330 -90436 80340 -89300
rect 80446 -90436 80456 -89300
rect 80508 -90436 80518 -89300
rect 80620 -90434 80630 -89298
rect 80682 -90434 80692 -89298
rect 80802 -90438 80812 -89302
rect 80864 -90438 80874 -89302
rect 80980 -90436 80990 -89300
rect 81042 -90436 81052 -89300
rect 81156 -90434 81166 -89298
rect 81218 -90434 81228 -89298
rect 81334 -90438 81344 -89302
rect 81396 -90438 81406 -89302
rect 81512 -90436 81522 -89300
rect 81574 -90436 81584 -89300
rect 81690 -90434 81700 -89298
rect 81752 -90434 81762 -89298
rect 81866 -90438 81876 -89302
rect 81928 -90438 81938 -89302
rect 82046 -90436 82056 -89300
rect 82108 -90436 82118 -89300
rect 82226 -90436 82236 -89300
rect 82288 -90436 82298 -89300
rect 82406 -90436 82416 -89300
rect 82468 -90436 82478 -89300
rect 82580 -90436 82590 -89300
rect 82642 -90436 82652 -89300
rect 82758 -90434 82768 -89298
rect 82820 -90434 82830 -89298
rect 82934 -90434 82944 -89298
rect 82996 -90434 83006 -89298
rect 83114 -90434 83124 -89298
rect 83176 -90434 83186 -89298
rect 83292 -90440 83302 -89304
rect 83354 -90440 83364 -89304
rect 83472 -90436 83482 -89300
rect 83534 -90436 83544 -89300
rect 83648 -90438 83658 -89302
rect 83710 -90438 83720 -89302
rect 83826 -90438 83836 -89302
rect 83888 -90438 83898 -89302
rect 84180 -91190 85972 -87756
rect 55044 -91892 55054 -91190
rect 85992 -91892 86002 -91190
<< via1 >>
rect 56256 -69858 64360 -69390
rect 68184 -69828 84246 -69294
rect 60954 -71284 61012 -70132
rect 61310 -71286 61368 -70134
rect 61664 -71286 61722 -70134
rect 62022 -71280 62080 -70128
rect 62376 -71286 62434 -70134
rect 62730 -71284 62788 -70132
rect 63090 -71282 63148 -70130
rect 63446 -71284 63504 -70132
rect 63802 -71282 63860 -70130
rect 64160 -71282 64218 -70130
rect 68128 -71254 68182 -70112
rect 68320 -71270 68374 -70128
rect 68488 -71270 68542 -70128
rect 68670 -71266 68724 -70124
rect 68848 -71262 68902 -70120
rect 69026 -71260 69080 -70118
rect 69200 -71262 69254 -70120
rect 69378 -71264 69432 -70122
rect 69558 -71262 69612 -70120
rect 69732 -71262 69786 -70120
rect 69910 -71262 69964 -70120
rect 70094 -71266 70148 -70124
rect 70268 -71262 70322 -70120
rect 70452 -71258 70506 -70116
rect 70620 -71262 70674 -70120
rect 70804 -71254 70858 -70112
rect 70980 -71256 71034 -70114
rect 71158 -71258 71212 -70116
rect 71336 -71256 71390 -70114
rect 71512 -71258 71566 -70116
rect 71694 -71258 71748 -70116
rect 71874 -71258 71928 -70116
rect 72046 -71262 72100 -70120
rect 72228 -71262 72282 -70120
rect 72406 -71262 72460 -70120
rect 72586 -71262 72640 -70120
rect 72756 -71262 72810 -70120
rect 72942 -71258 72996 -70116
rect 73122 -71258 73176 -70116
rect 73302 -71258 73356 -70116
rect 73472 -71264 73526 -70122
rect 73652 -71262 73706 -70120
rect 73832 -71258 73886 -70116
rect 74008 -71258 74062 -70116
rect 74180 -71256 74234 -70114
rect 74366 -71256 74420 -70114
rect 74540 -71258 74594 -70116
rect 74724 -71258 74778 -70116
rect 74896 -71258 74950 -70116
rect 75074 -71258 75128 -70116
rect 75252 -71256 75306 -70114
rect 75432 -71256 75486 -70114
rect 75610 -71258 75664 -70116
rect 75788 -71256 75842 -70114
rect 75966 -71254 76020 -70112
rect 76146 -71258 76200 -70116
rect 76320 -71258 76374 -70116
rect 76496 -71256 76550 -70114
rect 76674 -71258 76728 -70116
rect 76860 -71258 76914 -70116
rect 77036 -71258 77090 -70116
rect 77212 -71262 77266 -70120
rect 77392 -71258 77446 -70116
rect 77568 -71256 77622 -70114
rect 77744 -71262 77798 -70120
rect 77926 -71254 77980 -70112
rect 78104 -71258 78158 -70116
rect 78282 -71256 78336 -70114
rect 78452 -71258 78506 -70116
rect 78638 -71256 78692 -70114
rect 78812 -71262 78866 -70120
rect 78996 -71258 79050 -70116
rect 79170 -71258 79224 -70116
rect 79346 -71262 79400 -70120
rect 79522 -71258 79576 -70116
rect 79704 -71262 79758 -70120
rect 79882 -71262 79936 -70120
rect 80058 -71256 80112 -70114
rect 80236 -71258 80290 -70116
rect 80412 -71262 80466 -70120
rect 80594 -71262 80648 -70120
rect 80768 -71258 80822 -70116
rect 80948 -71256 81002 -70114
rect 81126 -71262 81180 -70120
rect 81306 -71258 81360 -70116
rect 81480 -71258 81534 -70116
rect 81660 -71262 81714 -70120
rect 81836 -71262 81890 -70120
rect 82010 -71262 82064 -70120
rect 82190 -71258 82244 -70116
rect 82374 -71258 82428 -70116
rect 82546 -71262 82600 -70120
rect 82726 -71258 82780 -70116
rect 82906 -71258 82960 -70116
rect 83086 -71258 83140 -70116
rect 83264 -71256 83318 -70114
rect 83440 -71264 83494 -70122
rect 83620 -71262 83674 -70120
rect 83796 -71262 83850 -70120
rect 83976 -71262 84030 -70120
rect 84154 -71264 84208 -70122
rect 68204 -71338 68302 -71328
rect 60846 -71343 60938 -71340
rect 61202 -71343 61294 -71342
rect 61558 -71343 61650 -71340
rect 61736 -71343 61828 -71340
rect 61916 -71343 62008 -71342
rect 62090 -71343 62182 -71342
rect 62448 -71343 62540 -71342
rect 62810 -71343 62902 -71342
rect 63338 -71343 63430 -71342
rect 63694 -71343 63786 -71342
rect 56330 -71484 59514 -71346
rect 60834 -71350 64295 -71343
rect 60834 -71406 64320 -71350
rect 60834 -71482 64295 -71406
rect 68200 -71482 68302 -71338
rect 68204 -71492 68302 -71482
rect 68374 -71482 68470 -71338
rect 68558 -71482 68654 -71338
rect 68734 -71482 68830 -71338
rect 68912 -71482 69008 -71338
rect 69092 -71482 69188 -71338
rect 69268 -71482 69364 -71338
rect 69444 -71480 69540 -71336
rect 69622 -71478 69718 -71334
rect 69800 -71480 69896 -71336
rect 69980 -71480 70076 -71336
rect 70158 -71482 70254 -71338
rect 70338 -71478 70434 -71334
rect 70514 -71482 70610 -71338
rect 70694 -71482 70790 -71338
rect 70874 -71480 70970 -71336
rect 71050 -71480 71146 -71336
rect 71228 -71482 71324 -71338
rect 71404 -71482 71500 -71338
rect 71580 -71480 71676 -71336
rect 71764 -71478 71860 -71334
rect 71940 -71482 72036 -71338
rect 72118 -71480 72214 -71336
rect 72294 -71480 72390 -71336
rect 72470 -71480 72566 -71336
rect 72648 -71478 72744 -71334
rect 72832 -71480 72928 -71336
rect 73006 -71480 73102 -71336
rect 73186 -71480 73282 -71336
rect 73362 -71482 73458 -71338
rect 73542 -71482 73638 -71338
rect 73720 -71482 73816 -71338
rect 73900 -71482 73996 -71338
rect 74074 -71480 74170 -71336
rect 74256 -71478 74352 -71334
rect 74434 -71480 74530 -71336
rect 74614 -71478 74710 -71334
rect 74792 -71476 74888 -71332
rect 74968 -71478 75064 -71334
rect 75146 -71480 75242 -71336
rect 75326 -71478 75422 -71334
rect 75502 -71482 75598 -71338
rect 75680 -71478 75776 -71334
rect 75856 -71478 75952 -71334
rect 76034 -71478 76130 -71334
rect 76214 -71478 76310 -71334
rect 76392 -71480 76488 -71336
rect 76572 -71478 76668 -71334
rect 76746 -71480 76842 -71336
rect 76922 -71480 77018 -71336
rect 77102 -71480 77198 -71336
rect 77282 -71480 77378 -71336
rect 77458 -71482 77554 -71338
rect 77636 -71480 77732 -71336
rect 77814 -71480 77910 -71336
rect 77990 -71478 78086 -71334
rect 78168 -71478 78264 -71334
rect 78348 -71478 78444 -71334
rect 78526 -71478 78622 -71334
rect 78704 -71478 78800 -71334
rect 78882 -71478 78978 -71334
rect 79062 -71478 79158 -71334
rect 79236 -71480 79332 -71336
rect 79412 -71482 79508 -71338
rect 79592 -71480 79688 -71336
rect 79770 -71480 79866 -71336
rect 79948 -71480 80044 -71336
rect 80126 -71480 80222 -71336
rect 80304 -71480 80400 -71336
rect 80484 -71480 80580 -71336
rect 80662 -71480 80758 -71336
rect 80840 -71478 80936 -71334
rect 81016 -71478 81112 -71334
rect 81198 -71478 81294 -71334
rect 81372 -71478 81468 -71334
rect 81554 -71478 81650 -71334
rect 81732 -71480 81828 -71336
rect 81908 -71480 82004 -71336
rect 82086 -71478 82182 -71334
rect 82264 -71478 82360 -71334
rect 82444 -71480 82540 -71336
rect 82622 -71480 82718 -71336
rect 82798 -71480 82894 -71336
rect 82980 -71480 83076 -71336
rect 83158 -71480 83254 -71336
rect 83334 -71478 83430 -71334
rect 83512 -71478 83608 -71334
rect 83688 -71478 83784 -71334
rect 83868 -71480 83964 -71336
rect 84046 -71480 84142 -71336
rect 68132 -72706 68190 -71562
rect 68314 -72706 68372 -71562
rect 68494 -72698 68552 -71554
rect 68668 -72698 68726 -71554
rect 68848 -72698 68906 -71554
rect 69028 -72698 69086 -71554
rect 69202 -72700 69260 -71556
rect 69382 -72702 69440 -71558
rect 69556 -72698 69614 -71554
rect 69740 -72706 69798 -71562
rect 69910 -72704 69968 -71560
rect 70092 -72704 70150 -71560
rect 70266 -72706 70324 -71562
rect 70444 -72704 70502 -71560
rect 70624 -72702 70682 -71558
rect 70800 -72704 70858 -71560
rect 70982 -72700 71040 -71556
rect 71156 -72702 71214 -71558
rect 71336 -72704 71394 -71560
rect 71516 -72702 71574 -71558
rect 71692 -72704 71750 -71560
rect 71870 -72702 71928 -71558
rect 72048 -72702 72106 -71558
rect 72230 -72702 72288 -71558
rect 72404 -72706 72462 -71562
rect 72586 -72704 72644 -71560
rect 72754 -72704 72812 -71560
rect 72938 -72702 72996 -71558
rect 73118 -72702 73176 -71558
rect 73292 -72706 73350 -71562
rect 73466 -72700 73524 -71556
rect 73654 -72704 73712 -71560
rect 73830 -72698 73888 -71554
rect 74010 -72698 74068 -71554
rect 74188 -72700 74246 -71556
rect 74364 -72696 74422 -71552
rect 74544 -72696 74602 -71552
rect 74720 -72698 74778 -71554
rect 74898 -72698 74956 -71554
rect 75078 -72708 75136 -71564
rect 75246 -72706 75304 -71562
rect 75432 -72702 75490 -71558
rect 75608 -72716 75666 -71572
rect 75786 -72708 75844 -71564
rect 75964 -72708 76022 -71564
rect 76146 -72700 76204 -71556
rect 76326 -72696 76384 -71552
rect 76500 -72700 76558 -71556
rect 76674 -72706 76732 -71562
rect 76854 -72706 76912 -71562
rect 77034 -72704 77092 -71560
rect 77212 -72706 77270 -71562
rect 77386 -72708 77444 -71564
rect 77566 -72706 77624 -71562
rect 77744 -72702 77802 -71558
rect 77924 -72708 77982 -71564
rect 78104 -72706 78162 -71562
rect 78276 -72712 78334 -71568
rect 78458 -72714 78516 -71570
rect 78636 -72712 78694 -71568
rect 78810 -72706 78868 -71562
rect 78990 -72712 79048 -71568
rect 79170 -72708 79228 -71564
rect 79344 -72710 79402 -71566
rect 79526 -72706 79584 -71562
rect 79700 -72706 79758 -71562
rect 79882 -72704 79940 -71560
rect 80058 -72704 80116 -71560
rect 80232 -72704 80290 -71560
rect 80416 -72702 80474 -71558
rect 80590 -72700 80648 -71556
rect 80772 -72706 80830 -71562
rect 80946 -72702 81004 -71558
rect 81124 -72704 81182 -71560
rect 81298 -72700 81356 -71556
rect 81482 -72700 81540 -71556
rect 81658 -72700 81716 -71556
rect 81836 -72700 81894 -71556
rect 82018 -72702 82076 -71558
rect 82196 -72704 82254 -71560
rect 82370 -72706 82428 -71562
rect 82556 -72702 82614 -71558
rect 82724 -72704 82782 -71560
rect 82908 -72698 82966 -71554
rect 83080 -72698 83138 -71554
rect 83262 -72698 83320 -71554
rect 83444 -72704 83502 -71560
rect 83622 -72706 83680 -71562
rect 83796 -72706 83854 -71562
rect 83978 -72700 84036 -71556
rect 84148 -72710 84206 -71566
rect 56314 -74544 56368 -73398
rect 56490 -74542 56544 -73396
rect 56668 -74546 56722 -73400
rect 56852 -74542 56906 -73396
rect 57026 -74550 57080 -73404
rect 57202 -74554 57256 -73408
rect 57382 -74550 57436 -73404
rect 57558 -74546 57612 -73400
rect 57740 -74546 57794 -73400
rect 57916 -74550 57970 -73404
rect 58094 -74550 58148 -73404
rect 58276 -74554 58330 -73408
rect 58450 -74550 58504 -73404
rect 58630 -74548 58684 -73402
rect 58806 -74548 58860 -73402
rect 58986 -74546 59040 -73400
rect 59166 -74546 59220 -73400
rect 59344 -74546 59398 -73400
rect 59522 -74542 59576 -73396
rect 59698 -74546 59752 -73400
rect 59876 -74550 59930 -73404
rect 60054 -74550 60108 -73404
rect 60228 -74550 60282 -73404
rect 60406 -74554 60460 -73408
rect 60588 -74554 60642 -73408
rect 60768 -74546 60822 -73400
rect 60944 -74550 60998 -73404
rect 61122 -74550 61176 -73404
rect 61298 -74554 61352 -73408
rect 61478 -74548 61532 -73402
rect 61656 -74546 61710 -73400
rect 61828 -74550 61882 -73404
rect 62008 -74550 62062 -73404
rect 62188 -74550 62242 -73404
rect 62368 -74550 62422 -73404
rect 62546 -74548 62600 -73402
rect 62720 -74544 62774 -73398
rect 62898 -74550 62952 -73404
rect 63080 -74548 63134 -73402
rect 63256 -74544 63310 -73398
rect 63432 -74548 63486 -73402
rect 63612 -74546 63666 -73400
rect 63790 -74546 63844 -73400
rect 63968 -74544 64022 -73398
rect 64146 -74542 64200 -73396
rect 64322 -74546 64376 -73400
rect 56364 -74792 56470 -74636
rect 56546 -74798 56652 -74642
rect 56728 -74794 56834 -74638
rect 56908 -74794 57014 -74638
rect 57086 -74792 57192 -74636
rect 57262 -74792 57368 -74636
rect 57446 -74794 57552 -74638
rect 57620 -74794 57726 -74638
rect 57794 -74794 57900 -74638
rect 57976 -74798 58082 -74642
rect 58150 -74794 58256 -74638
rect 58328 -74794 58434 -74638
rect 58508 -74794 58614 -74638
rect 58678 -74794 58784 -74638
rect 58858 -74794 58964 -74638
rect 59042 -74794 59148 -74638
rect 59216 -74794 59322 -74638
rect 59390 -74792 59496 -74636
rect 59568 -74788 59674 -74632
rect 59750 -74798 59856 -74642
rect 59926 -74794 60032 -74638
rect 60106 -74794 60212 -74638
rect 60278 -74794 60384 -74638
rect 60462 -74798 60568 -74642
rect 60636 -74794 60742 -74638
rect 60816 -74798 60922 -74642
rect 60992 -74798 61098 -74642
rect 61168 -74794 61274 -74638
rect 61348 -74798 61454 -74642
rect 61528 -74794 61634 -74638
rect 61706 -74802 61812 -74646
rect 61886 -74794 61992 -74638
rect 62062 -74798 62168 -74642
rect 62240 -74788 62346 -74632
rect 62418 -74794 62524 -74638
rect 62596 -74794 62702 -74638
rect 62776 -74798 62882 -74642
rect 62956 -74798 63062 -74642
rect 63130 -74794 63236 -74638
rect 63314 -74798 63420 -74642
rect 63482 -74798 63588 -74642
rect 63660 -74804 63766 -74648
rect 63848 -74792 63954 -74636
rect 64020 -74794 64126 -74638
rect 64200 -74792 64306 -74636
rect 56298 -76006 56352 -74860
rect 56474 -76004 56528 -74858
rect 56652 -76008 56706 -74862
rect 56836 -76004 56890 -74858
rect 57010 -76012 57064 -74866
rect 57186 -76016 57240 -74870
rect 57366 -76012 57420 -74866
rect 57542 -76008 57596 -74862
rect 57724 -76008 57778 -74862
rect 57900 -76012 57954 -74866
rect 58078 -76012 58132 -74866
rect 58260 -76016 58314 -74870
rect 58434 -76012 58488 -74866
rect 58614 -76010 58668 -74864
rect 58790 -76010 58844 -74864
rect 58970 -76008 59024 -74862
rect 59150 -76008 59204 -74862
rect 59328 -76008 59382 -74862
rect 59506 -76004 59560 -74858
rect 59682 -76008 59736 -74862
rect 59860 -76012 59914 -74866
rect 60038 -76012 60092 -74866
rect 60212 -76012 60266 -74866
rect 60390 -76016 60444 -74870
rect 60572 -76016 60626 -74870
rect 60752 -76008 60806 -74862
rect 60928 -76012 60982 -74866
rect 61106 -76012 61160 -74866
rect 61282 -76016 61336 -74870
rect 61462 -76010 61516 -74864
rect 61640 -76008 61694 -74862
rect 61812 -76012 61866 -74866
rect 61992 -76012 62046 -74866
rect 62172 -76012 62226 -74866
rect 62352 -76012 62406 -74866
rect 62530 -76010 62584 -74864
rect 62704 -76006 62758 -74860
rect 62882 -76012 62936 -74866
rect 63064 -76010 63118 -74864
rect 63240 -76006 63294 -74860
rect 63416 -76010 63470 -74864
rect 63596 -76008 63650 -74862
rect 63774 -76008 63828 -74862
rect 63952 -76006 64006 -74860
rect 64130 -76004 64184 -74858
rect 64306 -76008 64360 -74862
rect 56304 -78394 56358 -77248
rect 56480 -78392 56534 -77246
rect 56658 -78396 56712 -77250
rect 56842 -78392 56896 -77246
rect 57016 -78400 57070 -77254
rect 57192 -78404 57246 -77258
rect 57372 -78400 57426 -77254
rect 57548 -78396 57602 -77250
rect 57730 -78396 57784 -77250
rect 57906 -78400 57960 -77254
rect 58084 -78400 58138 -77254
rect 58266 -78404 58320 -77258
rect 58440 -78400 58494 -77254
rect 58620 -78398 58674 -77252
rect 58796 -78398 58850 -77252
rect 58976 -78396 59030 -77250
rect 59156 -78396 59210 -77250
rect 59334 -78396 59388 -77250
rect 59512 -78392 59566 -77246
rect 59688 -78396 59742 -77250
rect 59866 -78400 59920 -77254
rect 60044 -78400 60098 -77254
rect 60218 -78400 60272 -77254
rect 60396 -78404 60450 -77258
rect 60578 -78404 60632 -77258
rect 60758 -78396 60812 -77250
rect 60934 -78400 60988 -77254
rect 61112 -78400 61166 -77254
rect 61288 -78404 61342 -77258
rect 61468 -78398 61522 -77252
rect 61646 -78396 61700 -77250
rect 61818 -78400 61872 -77254
rect 61998 -78400 62052 -77254
rect 62178 -78400 62232 -77254
rect 62358 -78400 62412 -77254
rect 62536 -78398 62590 -77252
rect 62710 -78394 62764 -77248
rect 62888 -78400 62942 -77254
rect 63070 -78398 63124 -77252
rect 63246 -78394 63300 -77248
rect 63422 -78398 63476 -77252
rect 63602 -78396 63656 -77250
rect 63780 -78396 63834 -77250
rect 63958 -78394 64012 -77248
rect 64136 -78392 64190 -77246
rect 64312 -78396 64366 -77250
rect 56354 -78642 56460 -78486
rect 56536 -78648 56642 -78492
rect 56718 -78644 56824 -78488
rect 56898 -78644 57004 -78488
rect 57076 -78642 57182 -78486
rect 57252 -78642 57358 -78486
rect 57436 -78644 57542 -78488
rect 57610 -78644 57716 -78488
rect 57784 -78644 57890 -78488
rect 57966 -78648 58072 -78492
rect 58140 -78644 58246 -78488
rect 58318 -78644 58424 -78488
rect 58498 -78644 58604 -78488
rect 58668 -78644 58774 -78488
rect 58848 -78644 58954 -78488
rect 59032 -78644 59138 -78488
rect 59206 -78644 59312 -78488
rect 59380 -78642 59486 -78486
rect 59558 -78638 59664 -78482
rect 59740 -78648 59846 -78492
rect 59916 -78644 60022 -78488
rect 60096 -78644 60202 -78488
rect 60268 -78644 60374 -78488
rect 60452 -78648 60558 -78492
rect 60626 -78644 60732 -78488
rect 60806 -78648 60912 -78492
rect 60982 -78648 61088 -78492
rect 61158 -78644 61264 -78488
rect 61338 -78648 61444 -78492
rect 61518 -78644 61624 -78488
rect 61696 -78652 61802 -78496
rect 61876 -78644 61982 -78488
rect 62052 -78648 62158 -78492
rect 62230 -78638 62336 -78482
rect 62408 -78644 62514 -78488
rect 62586 -78644 62692 -78488
rect 62766 -78648 62872 -78492
rect 62946 -78648 63052 -78492
rect 63120 -78644 63226 -78488
rect 63304 -78648 63410 -78492
rect 63472 -78648 63578 -78492
rect 63650 -78654 63756 -78498
rect 63838 -78642 63944 -78486
rect 64010 -78644 64116 -78488
rect 64190 -78642 64296 -78486
rect 56288 -79856 56342 -78710
rect 56464 -79854 56518 -78708
rect 56642 -79858 56696 -78712
rect 56826 -79854 56880 -78708
rect 57000 -79862 57054 -78716
rect 57176 -79866 57230 -78720
rect 57356 -79862 57410 -78716
rect 57532 -79858 57586 -78712
rect 57714 -79858 57768 -78712
rect 57890 -79862 57944 -78716
rect 58068 -79862 58122 -78716
rect 58250 -79866 58304 -78720
rect 58424 -79862 58478 -78716
rect 58604 -79860 58658 -78714
rect 58780 -79860 58834 -78714
rect 58960 -79858 59014 -78712
rect 59140 -79858 59194 -78712
rect 59318 -79858 59372 -78712
rect 59496 -79854 59550 -78708
rect 59672 -79858 59726 -78712
rect 59850 -79862 59904 -78716
rect 60028 -79862 60082 -78716
rect 60202 -79862 60256 -78716
rect 60380 -79866 60434 -78720
rect 60562 -79866 60616 -78720
rect 60742 -79858 60796 -78712
rect 60918 -79862 60972 -78716
rect 61096 -79862 61150 -78716
rect 61272 -79866 61326 -78720
rect 61452 -79860 61506 -78714
rect 61630 -79858 61684 -78712
rect 61802 -79862 61856 -78716
rect 61982 -79862 62036 -78716
rect 62162 -79862 62216 -78716
rect 62342 -79862 62396 -78716
rect 62520 -79860 62574 -78714
rect 62694 -79856 62748 -78710
rect 62872 -79862 62926 -78716
rect 63054 -79860 63108 -78714
rect 63230 -79856 63284 -78710
rect 63406 -79860 63460 -78714
rect 63586 -79858 63640 -78712
rect 63764 -79858 63818 -78712
rect 63942 -79856 63996 -78710
rect 64120 -79854 64174 -78708
rect 64296 -79858 64350 -78712
rect 56314 -82360 56368 -81214
rect 56490 -82358 56544 -81212
rect 56668 -82362 56722 -81216
rect 56852 -82358 56906 -81212
rect 57026 -82366 57080 -81220
rect 57202 -82370 57256 -81224
rect 57382 -82366 57436 -81220
rect 57558 -82362 57612 -81216
rect 57740 -82362 57794 -81216
rect 57916 -82366 57970 -81220
rect 58094 -82366 58148 -81220
rect 58276 -82370 58330 -81224
rect 58450 -82366 58504 -81220
rect 58630 -82364 58684 -81218
rect 58806 -82364 58860 -81218
rect 58986 -82362 59040 -81216
rect 59166 -82362 59220 -81216
rect 59344 -82362 59398 -81216
rect 59522 -82358 59576 -81212
rect 59698 -82362 59752 -81216
rect 59876 -82366 59930 -81220
rect 60054 -82366 60108 -81220
rect 60228 -82366 60282 -81220
rect 60406 -82370 60460 -81224
rect 60588 -82370 60642 -81224
rect 60768 -82362 60822 -81216
rect 60944 -82366 60998 -81220
rect 61122 -82366 61176 -81220
rect 61298 -82370 61352 -81224
rect 61478 -82364 61532 -81218
rect 61656 -82362 61710 -81216
rect 61828 -82366 61882 -81220
rect 62008 -82366 62062 -81220
rect 62188 -82366 62242 -81220
rect 62368 -82366 62422 -81220
rect 62546 -82364 62600 -81218
rect 62720 -82360 62774 -81214
rect 62898 -82366 62952 -81220
rect 63080 -82364 63134 -81218
rect 63256 -82360 63310 -81214
rect 63432 -82364 63486 -81218
rect 63612 -82362 63666 -81216
rect 63790 -82362 63844 -81216
rect 63968 -82360 64022 -81214
rect 64146 -82358 64200 -81212
rect 64322 -82362 64376 -81216
rect 56364 -82608 56470 -82452
rect 56546 -82614 56652 -82458
rect 56728 -82610 56834 -82454
rect 56908 -82610 57014 -82454
rect 57086 -82608 57192 -82452
rect 57262 -82608 57368 -82452
rect 57446 -82610 57552 -82454
rect 57620 -82610 57726 -82454
rect 57794 -82610 57900 -82454
rect 57976 -82614 58082 -82458
rect 58150 -82610 58256 -82454
rect 58328 -82610 58434 -82454
rect 58508 -82610 58614 -82454
rect 58678 -82610 58784 -82454
rect 58858 -82610 58964 -82454
rect 59042 -82610 59148 -82454
rect 59216 -82610 59322 -82454
rect 59390 -82608 59496 -82452
rect 59568 -82604 59674 -82448
rect 59750 -82614 59856 -82458
rect 59926 -82610 60032 -82454
rect 60106 -82610 60212 -82454
rect 60278 -82610 60384 -82454
rect 60462 -82614 60568 -82458
rect 60636 -82610 60742 -82454
rect 60816 -82614 60922 -82458
rect 60992 -82614 61098 -82458
rect 61168 -82610 61274 -82454
rect 61348 -82614 61454 -82458
rect 61528 -82610 61634 -82454
rect 61706 -82618 61812 -82462
rect 61886 -82610 61992 -82454
rect 62062 -82614 62168 -82458
rect 62240 -82604 62346 -82448
rect 62418 -82610 62524 -82454
rect 62596 -82610 62702 -82454
rect 62776 -82614 62882 -82458
rect 62956 -82614 63062 -82458
rect 63130 -82610 63236 -82454
rect 63314 -82614 63420 -82458
rect 63482 -82614 63588 -82458
rect 63660 -82620 63766 -82464
rect 63848 -82608 63954 -82452
rect 64020 -82610 64126 -82454
rect 64200 -82608 64306 -82452
rect 56298 -83822 56352 -82676
rect 56474 -83820 56528 -82674
rect 56652 -83824 56706 -82678
rect 56836 -83820 56890 -82674
rect 57010 -83828 57064 -82682
rect 57186 -83832 57240 -82686
rect 57366 -83828 57420 -82682
rect 57542 -83824 57596 -82678
rect 57724 -83824 57778 -82678
rect 57900 -83828 57954 -82682
rect 58078 -83828 58132 -82682
rect 58260 -83832 58314 -82686
rect 58434 -83828 58488 -82682
rect 58614 -83826 58668 -82680
rect 58790 -83826 58844 -82680
rect 58970 -83824 59024 -82678
rect 59150 -83824 59204 -82678
rect 59328 -83824 59382 -82678
rect 59506 -83820 59560 -82674
rect 59682 -83824 59736 -82678
rect 59860 -83828 59914 -82682
rect 60038 -83828 60092 -82682
rect 60212 -83828 60266 -82682
rect 60390 -83832 60444 -82686
rect 60572 -83832 60626 -82686
rect 60752 -83824 60806 -82678
rect 60928 -83828 60982 -82682
rect 61106 -83828 61160 -82682
rect 61282 -83832 61336 -82686
rect 61462 -83826 61516 -82680
rect 61640 -83824 61694 -82678
rect 61812 -83828 61866 -82682
rect 61992 -83828 62046 -82682
rect 62172 -83828 62226 -82682
rect 62352 -83828 62406 -82682
rect 62530 -83826 62584 -82680
rect 62704 -83822 62758 -82676
rect 62882 -83828 62936 -82682
rect 63064 -83826 63118 -82680
rect 63240 -83822 63294 -82676
rect 63416 -83826 63470 -82680
rect 63596 -83824 63650 -82678
rect 63774 -83824 63828 -82678
rect 63952 -83822 64006 -82676
rect 64130 -83820 64184 -82674
rect 64306 -83824 64360 -82678
rect 56286 -86180 56340 -85034
rect 56462 -86178 56516 -85032
rect 56640 -86182 56694 -85036
rect 56824 -86178 56878 -85032
rect 56998 -86186 57052 -85040
rect 57174 -86190 57228 -85044
rect 57354 -86186 57408 -85040
rect 57530 -86182 57584 -85036
rect 57712 -86182 57766 -85036
rect 57888 -86186 57942 -85040
rect 58066 -86186 58120 -85040
rect 58248 -86190 58302 -85044
rect 58422 -86186 58476 -85040
rect 58602 -86184 58656 -85038
rect 58778 -86184 58832 -85038
rect 58958 -86182 59012 -85036
rect 59138 -86182 59192 -85036
rect 59316 -86182 59370 -85036
rect 59494 -86178 59548 -85032
rect 59670 -86182 59724 -85036
rect 59848 -86186 59902 -85040
rect 60026 -86186 60080 -85040
rect 60200 -86186 60254 -85040
rect 60378 -86190 60432 -85044
rect 60560 -86190 60614 -85044
rect 60740 -86182 60794 -85036
rect 60916 -86186 60970 -85040
rect 61094 -86186 61148 -85040
rect 61270 -86190 61324 -85044
rect 61450 -86184 61504 -85038
rect 61628 -86182 61682 -85036
rect 61800 -86186 61854 -85040
rect 61980 -86186 62034 -85040
rect 62160 -86186 62214 -85040
rect 62340 -86186 62394 -85040
rect 62518 -86184 62572 -85038
rect 62692 -86180 62746 -85034
rect 62870 -86186 62924 -85040
rect 63052 -86184 63106 -85038
rect 63228 -86180 63282 -85034
rect 63404 -86184 63458 -85038
rect 63584 -86182 63638 -85036
rect 63762 -86182 63816 -85036
rect 63940 -86180 63994 -85034
rect 64118 -86178 64172 -85032
rect 64294 -86182 64348 -85036
rect 56336 -86428 56442 -86272
rect 56518 -86434 56624 -86278
rect 56700 -86430 56806 -86274
rect 56880 -86430 56986 -86274
rect 57058 -86428 57164 -86272
rect 57234 -86428 57340 -86272
rect 57418 -86430 57524 -86274
rect 57592 -86430 57698 -86274
rect 57766 -86430 57872 -86274
rect 57948 -86434 58054 -86278
rect 58122 -86430 58228 -86274
rect 58300 -86430 58406 -86274
rect 58480 -86430 58586 -86274
rect 58650 -86430 58756 -86274
rect 58830 -86430 58936 -86274
rect 59014 -86430 59120 -86274
rect 59188 -86430 59294 -86274
rect 59362 -86428 59468 -86272
rect 59540 -86424 59646 -86268
rect 59722 -86434 59828 -86278
rect 59898 -86430 60004 -86274
rect 60078 -86430 60184 -86274
rect 60250 -86430 60356 -86274
rect 60434 -86434 60540 -86278
rect 60608 -86430 60714 -86274
rect 60788 -86434 60894 -86278
rect 60964 -86434 61070 -86278
rect 61140 -86430 61246 -86274
rect 61320 -86434 61426 -86278
rect 61500 -86430 61606 -86274
rect 61678 -86438 61784 -86282
rect 61858 -86430 61964 -86274
rect 62034 -86434 62140 -86278
rect 62212 -86424 62318 -86268
rect 62390 -86430 62496 -86274
rect 62568 -86430 62674 -86274
rect 62748 -86434 62854 -86278
rect 62928 -86434 63034 -86278
rect 63102 -86430 63208 -86274
rect 63286 -86434 63392 -86278
rect 63454 -86434 63560 -86278
rect 63632 -86440 63738 -86284
rect 63820 -86428 63926 -86272
rect 63992 -86430 64098 -86274
rect 64172 -86428 64278 -86272
rect 56270 -87642 56324 -86496
rect 56446 -87640 56500 -86494
rect 56624 -87644 56678 -86498
rect 56808 -87640 56862 -86494
rect 56982 -87648 57036 -86502
rect 57158 -87652 57212 -86506
rect 57338 -87648 57392 -86502
rect 57514 -87644 57568 -86498
rect 57696 -87644 57750 -86498
rect 57872 -87648 57926 -86502
rect 58050 -87648 58104 -86502
rect 58232 -87652 58286 -86506
rect 58406 -87648 58460 -86502
rect 58586 -87646 58640 -86500
rect 58762 -87646 58816 -86500
rect 58942 -87644 58996 -86498
rect 59122 -87644 59176 -86498
rect 59300 -87644 59354 -86498
rect 59478 -87640 59532 -86494
rect 59654 -87644 59708 -86498
rect 59832 -87648 59886 -86502
rect 60010 -87648 60064 -86502
rect 60184 -87648 60238 -86502
rect 60362 -87652 60416 -86506
rect 60544 -87652 60598 -86506
rect 60724 -87644 60778 -86498
rect 60900 -87648 60954 -86502
rect 61078 -87648 61132 -86502
rect 61254 -87652 61308 -86506
rect 61434 -87646 61488 -86500
rect 61612 -87644 61666 -86498
rect 61784 -87648 61838 -86502
rect 61964 -87648 62018 -86502
rect 62144 -87648 62198 -86502
rect 62324 -87648 62378 -86502
rect 62502 -87646 62556 -86500
rect 62676 -87642 62730 -86496
rect 62854 -87648 62908 -86502
rect 63036 -87646 63090 -86500
rect 63212 -87642 63266 -86496
rect 63388 -87646 63442 -86500
rect 63568 -87644 63622 -86498
rect 63746 -87644 63800 -86498
rect 63924 -87642 63978 -86496
rect 64102 -87640 64156 -86494
rect 64278 -87644 64332 -86498
rect 66140 -87790 66196 -87616
rect 66318 -87788 66374 -87614
rect 66498 -87786 66554 -87612
rect 66676 -87788 66732 -87614
rect 66848 -87788 66904 -87614
rect 67030 -87786 67086 -87612
rect 67208 -87786 67264 -87612
rect 55742 -88354 56040 -87954
rect 66212 -87990 66316 -87838
rect 66392 -87990 66496 -87838
rect 66570 -87990 66674 -87838
rect 66746 -87990 66850 -87838
rect 66924 -87990 67028 -87838
rect 67100 -87990 67204 -87838
rect 66146 -88218 66202 -88044
rect 66326 -88214 66382 -88040
rect 66506 -88216 66562 -88042
rect 66684 -88216 66740 -88042
rect 66862 -88216 66918 -88042
rect 67040 -88216 67096 -88042
rect 67218 -88220 67274 -88046
rect 66136 -88626 66192 -88452
rect 66320 -88620 66376 -88446
rect 66500 -88624 66556 -88450
rect 66676 -88626 66732 -88452
rect 66854 -88620 66910 -88446
rect 67034 -88622 67090 -88448
rect 67212 -88626 67268 -88452
rect 66210 -88826 66314 -88674
rect 66392 -88828 66496 -88676
rect 66564 -88830 66668 -88678
rect 66746 -88830 66850 -88678
rect 66924 -88830 67028 -88678
rect 67104 -88830 67208 -88678
rect 66140 -89028 66192 -88874
rect 66320 -89034 66372 -88880
rect 66496 -89030 66548 -88876
rect 66672 -89034 66724 -88880
rect 66852 -89036 66904 -88882
rect 67034 -89034 67086 -88880
rect 67224 -89036 67276 -88882
rect 68260 -89018 68312 -87882
rect 68442 -89012 68494 -87876
rect 68628 -89020 68680 -87884
rect 68802 -89026 68854 -87890
rect 68980 -89026 69032 -87890
rect 69160 -89026 69212 -87890
rect 69336 -89026 69388 -87890
rect 69514 -89022 69566 -87886
rect 69694 -89024 69746 -87888
rect 69868 -89022 69920 -87886
rect 70048 -89026 70100 -87890
rect 70224 -89024 70276 -87888
rect 70404 -89024 70456 -87888
rect 70582 -89026 70634 -87890
rect 70760 -89028 70812 -87892
rect 70936 -89026 70988 -87890
rect 71114 -89028 71166 -87892
rect 71294 -89026 71346 -87890
rect 71472 -89026 71524 -87890
rect 71648 -89028 71700 -87892
rect 71826 -89026 71878 -87890
rect 56418 -89246 56534 -89192
rect 56598 -89248 56714 -89194
rect 56784 -89248 56900 -89194
rect 56968 -89246 57084 -89192
rect 57144 -89246 57260 -89192
rect 57318 -89246 57434 -89192
rect 57494 -89248 57610 -89194
rect 57682 -89254 57798 -89200
rect 57856 -89254 57972 -89200
rect 58038 -89266 58154 -89212
rect 58214 -89268 58292 -89210
rect 58412 -89266 58490 -89208
rect 58574 -89266 58652 -89208
rect 58760 -89266 58838 -89208
rect 58936 -89268 59014 -89210
rect 59108 -89266 59186 -89208
rect 59292 -89266 59370 -89208
rect 59468 -89262 59546 -89204
rect 59642 -89262 59720 -89204
rect 59832 -89266 59910 -89208
rect 60874 -89262 60952 -89204
rect 61064 -89266 61142 -89208
rect 61242 -89268 61320 -89210
rect 61416 -89262 61494 -89204
rect 61594 -89254 61672 -89196
rect 61770 -89262 61848 -89204
rect 61962 -89262 62040 -89204
rect 62122 -89258 62200 -89200
rect 62298 -89262 62376 -89204
rect 62478 -89262 62556 -89204
rect 62652 -89266 62730 -89208
rect 62842 -89258 62920 -89200
rect 63026 -89258 63104 -89200
rect 63188 -89258 63266 -89200
rect 63370 -89262 63448 -89204
rect 63554 -89266 63632 -89208
rect 63716 -89258 63794 -89200
rect 63900 -89258 63978 -89200
rect 64088 -89258 64166 -89200
rect 64256 -89258 64334 -89200
rect 56362 -90484 56414 -89326
rect 56548 -90484 56600 -89326
rect 56720 -90492 56772 -89334
rect 56906 -90484 56958 -89326
rect 57072 -90484 57124 -89326
rect 57260 -90484 57312 -89326
rect 57434 -90486 57486 -89328
rect 57614 -90486 57666 -89328
rect 57780 -90486 57832 -89328
rect 57974 -90484 58026 -89326
rect 58142 -90476 58194 -89318
rect 58328 -90480 58380 -89322
rect 58500 -90484 58552 -89326
rect 58686 -90480 58738 -89322
rect 58858 -90484 58910 -89326
rect 59038 -90486 59090 -89328
rect 59214 -90488 59266 -89330
rect 59396 -90486 59448 -89328
rect 59570 -90484 59622 -89326
rect 59752 -90484 59804 -89326
rect 59922 -90480 59974 -89322
rect 60796 -90484 60848 -89326
rect 60980 -90484 61032 -89326
rect 61142 -90484 61194 -89326
rect 61330 -90486 61382 -89328
rect 61506 -90486 61558 -89328
rect 61690 -90486 61742 -89328
rect 61862 -90490 61914 -89332
rect 62042 -90484 62094 -89326
rect 62216 -90480 62268 -89322
rect 62398 -90484 62450 -89326
rect 62570 -90480 62622 -89322
rect 62756 -90484 62808 -89326
rect 62926 -90484 62978 -89326
rect 63112 -90478 63164 -89320
rect 63288 -90480 63340 -89322
rect 63468 -90486 63520 -89328
rect 63638 -90490 63690 -89332
rect 63826 -90484 63878 -89326
rect 63994 -90486 64046 -89328
rect 64184 -90484 64236 -89326
rect 64348 -90486 64400 -89328
rect 68330 -89228 68424 -89082
rect 68510 -89228 68604 -89082
rect 68690 -89228 68784 -89082
rect 68868 -89228 68962 -89082
rect 69044 -89228 69138 -89082
rect 69224 -89230 69318 -89084
rect 69400 -89228 69494 -89082
rect 69578 -89228 69672 -89082
rect 69760 -89228 69854 -89082
rect 69934 -89226 70028 -89080
rect 70114 -89228 70208 -89082
rect 70290 -89230 70384 -89084
rect 70470 -89228 70564 -89082
rect 70644 -89226 70738 -89080
rect 70824 -89224 70918 -89078
rect 71002 -89228 71096 -89082
rect 71180 -89226 71274 -89080
rect 71360 -89228 71454 -89082
rect 71536 -89228 71630 -89082
rect 71714 -89228 71808 -89082
rect 68268 -90444 68320 -89308
rect 68446 -90444 68498 -89308
rect 68620 -90442 68672 -89306
rect 68802 -90446 68854 -89310
rect 68980 -90444 69032 -89308
rect 69156 -90442 69208 -89306
rect 69334 -90446 69386 -89310
rect 69512 -90444 69564 -89308
rect 69690 -90442 69742 -89306
rect 69866 -90446 69918 -89310
rect 70046 -90444 70098 -89308
rect 70226 -90444 70278 -89308
rect 70406 -90444 70458 -89308
rect 70580 -90444 70632 -89308
rect 70758 -90442 70810 -89306
rect 70934 -90442 70986 -89306
rect 71114 -90442 71166 -89306
rect 71292 -90448 71344 -89312
rect 71472 -90444 71524 -89308
rect 71648 -90446 71700 -89310
rect 71826 -90446 71878 -89310
rect 74156 -89016 74208 -87880
rect 74338 -89010 74390 -87874
rect 74524 -89018 74576 -87882
rect 74698 -89024 74750 -87888
rect 74876 -89024 74928 -87888
rect 75056 -89024 75108 -87888
rect 75232 -89024 75284 -87888
rect 75410 -89020 75462 -87884
rect 75590 -89022 75642 -87886
rect 75764 -89020 75816 -87884
rect 75944 -89024 75996 -87888
rect 76120 -89022 76172 -87886
rect 76300 -89022 76352 -87886
rect 76478 -89024 76530 -87888
rect 76656 -89026 76708 -87890
rect 76832 -89024 76884 -87888
rect 77010 -89026 77062 -87890
rect 77190 -89024 77242 -87888
rect 77368 -89024 77420 -87888
rect 77544 -89026 77596 -87890
rect 77722 -89024 77774 -87888
rect 74226 -89226 74320 -89080
rect 74406 -89226 74500 -89080
rect 74586 -89226 74680 -89080
rect 74764 -89226 74858 -89080
rect 74940 -89226 75034 -89080
rect 75120 -89228 75214 -89082
rect 75296 -89226 75390 -89080
rect 75474 -89226 75568 -89080
rect 75656 -89226 75750 -89080
rect 75830 -89224 75924 -89078
rect 76010 -89226 76104 -89080
rect 76186 -89228 76280 -89082
rect 76366 -89226 76460 -89080
rect 76540 -89224 76634 -89078
rect 76720 -89222 76814 -89076
rect 76898 -89226 76992 -89080
rect 77076 -89224 77170 -89078
rect 77256 -89226 77350 -89080
rect 77432 -89226 77526 -89080
rect 77610 -89226 77704 -89080
rect 74164 -90442 74216 -89306
rect 74342 -90442 74394 -89306
rect 74516 -90440 74568 -89304
rect 74698 -90444 74750 -89308
rect 74876 -90442 74928 -89306
rect 75052 -90440 75104 -89304
rect 75230 -90444 75282 -89308
rect 75408 -90442 75460 -89306
rect 75586 -90440 75638 -89304
rect 75762 -90444 75814 -89308
rect 75942 -90442 75994 -89306
rect 76122 -90442 76174 -89306
rect 76302 -90442 76354 -89306
rect 76476 -90442 76528 -89306
rect 76654 -90440 76706 -89304
rect 76830 -90440 76882 -89304
rect 77010 -90440 77062 -89304
rect 77188 -90446 77240 -89310
rect 77368 -90442 77420 -89306
rect 77544 -90444 77596 -89308
rect 77722 -90444 77774 -89308
rect 80270 -89010 80322 -87874
rect 80452 -89004 80504 -87868
rect 80638 -89012 80690 -87876
rect 80812 -89018 80864 -87882
rect 80990 -89018 81042 -87882
rect 81170 -89018 81222 -87882
rect 81346 -89018 81398 -87882
rect 81524 -89014 81576 -87878
rect 81704 -89016 81756 -87880
rect 81878 -89014 81930 -87878
rect 82058 -89018 82110 -87882
rect 82234 -89016 82286 -87880
rect 82414 -89016 82466 -87880
rect 82592 -89018 82644 -87882
rect 82770 -89020 82822 -87884
rect 82946 -89018 82998 -87882
rect 83124 -89020 83176 -87884
rect 83304 -89018 83356 -87882
rect 83482 -89018 83534 -87882
rect 83658 -89020 83710 -87884
rect 83836 -89018 83888 -87882
rect 80340 -89220 80434 -89074
rect 80520 -89220 80614 -89074
rect 80700 -89220 80794 -89074
rect 80878 -89220 80972 -89074
rect 81054 -89220 81148 -89074
rect 81234 -89222 81328 -89076
rect 81410 -89220 81504 -89074
rect 81588 -89220 81682 -89074
rect 81770 -89220 81864 -89074
rect 81944 -89218 82038 -89072
rect 82124 -89220 82218 -89074
rect 82300 -89222 82394 -89076
rect 82480 -89220 82574 -89074
rect 82654 -89218 82748 -89072
rect 82834 -89216 82928 -89070
rect 83012 -89220 83106 -89074
rect 83190 -89218 83284 -89072
rect 83370 -89220 83464 -89074
rect 83546 -89220 83640 -89074
rect 83724 -89220 83818 -89074
rect 80278 -90436 80330 -89300
rect 80456 -90436 80508 -89300
rect 80630 -90434 80682 -89298
rect 80812 -90438 80864 -89302
rect 80990 -90436 81042 -89300
rect 81166 -90434 81218 -89298
rect 81344 -90438 81396 -89302
rect 81522 -90436 81574 -89300
rect 81700 -90434 81752 -89298
rect 81876 -90438 81928 -89302
rect 82056 -90436 82108 -89300
rect 82236 -90436 82288 -89300
rect 82416 -90436 82468 -89300
rect 82590 -90436 82642 -89300
rect 82768 -90434 82820 -89298
rect 82944 -90434 82996 -89298
rect 83124 -90434 83176 -89298
rect 83302 -90440 83354 -89304
rect 83482 -90436 83534 -89300
rect 83658 -90438 83710 -89302
rect 83836 -90438 83888 -89302
rect 55054 -91892 85992 -91190
<< metal2 >>
rect 52320 -69294 86894 -69270
rect 52320 -69390 68184 -69294
rect 52320 -69842 56256 -69390
rect 64360 -69828 68184 -69390
rect 84246 -69828 86894 -69294
rect 64360 -69842 86894 -69828
rect 56256 -69868 64360 -69858
rect 68138 -70102 68180 -69842
rect 56462 -71336 56504 -70111
rect 56816 -71336 56858 -70107
rect 57182 -71336 57224 -70111
rect 57528 -71336 57570 -70111
rect 57892 -71336 57934 -70111
rect 58248 -71336 58290 -70107
rect 58604 -71336 58646 -70111
rect 58954 -71336 58996 -70107
rect 59312 -71336 59354 -70107
rect 68128 -70112 68182 -70102
rect 60962 -70122 60996 -70116
rect 60954 -70124 61012 -70122
rect 61318 -70124 61352 -70116
rect 61672 -70124 61706 -70116
rect 62030 -70118 62064 -70114
rect 62022 -70120 62080 -70118
rect 60946 -70132 61016 -70124
rect 61310 -70128 61368 -70124
rect 60946 -70134 60954 -70132
rect 61012 -70134 61016 -70132
rect 60946 -71294 61016 -71284
rect 61302 -70134 61372 -70128
rect 61664 -70132 61722 -70124
rect 62004 -70128 62080 -70120
rect 62386 -70124 62420 -70116
rect 62740 -70122 62774 -70114
rect 63096 -70120 63130 -70114
rect 63456 -70120 63490 -70114
rect 63812 -70118 63846 -70114
rect 62004 -70130 62022 -70128
rect 61302 -70138 61310 -70134
rect 61368 -70138 61372 -70134
rect 61302 -71298 61372 -71288
rect 61654 -70134 61724 -70132
rect 61654 -70142 61664 -70134
rect 61722 -70142 61724 -70134
rect 62376 -70134 62434 -70124
rect 62730 -70132 62788 -70122
rect 63088 -70130 63158 -70120
rect 62004 -71290 62080 -71280
rect 62366 -70144 62376 -70134
rect 62434 -70144 62436 -70134
rect 62030 -71292 62064 -71290
rect 61654 -71302 61724 -71292
rect 62366 -71304 62436 -71294
rect 62726 -70142 62730 -70132
rect 62788 -70142 62796 -70132
rect 63088 -71282 63090 -71280
rect 63148 -71282 63158 -71280
rect 63088 -71290 63158 -71282
rect 63436 -70130 63506 -70120
rect 63436 -71284 63446 -71280
rect 63504 -71284 63506 -71280
rect 63436 -71290 63506 -71284
rect 63794 -70128 63864 -70118
rect 63794 -71282 63802 -71278
rect 63860 -71282 63864 -71278
rect 63794 -71288 63864 -71282
rect 64150 -70124 64220 -70114
rect 68324 -70116 68358 -70094
rect 68128 -71264 68182 -71254
rect 68320 -70126 68382 -70116
rect 68490 -70118 68532 -69842
rect 68680 -70112 68714 -70094
rect 68854 -70110 68896 -69842
rect 69036 -70106 69070 -70094
rect 64150 -71282 64160 -71274
rect 64218 -71282 64220 -71274
rect 68138 -71279 68180 -71264
rect 68320 -71280 68382 -71270
rect 68488 -70128 68542 -70118
rect 68488 -71280 68542 -71270
rect 68670 -70122 68732 -70112
rect 68670 -71276 68732 -71266
rect 68848 -70120 68902 -70110
rect 68848 -71272 68902 -71262
rect 69026 -70116 69088 -70106
rect 69202 -70110 69244 -69842
rect 69392 -70110 69426 -70094
rect 69560 -70110 69602 -69842
rect 69748 -70108 69782 -70094
rect 69026 -71270 69088 -71260
rect 69200 -70120 69254 -70110
rect 69200 -71272 69254 -71262
rect 69378 -70120 69440 -70110
rect 64150 -71284 64220 -71282
rect 63090 -71292 63148 -71290
rect 62726 -71302 62796 -71292
rect 63446 -71294 63504 -71290
rect 63802 -71292 63860 -71288
rect 64160 -71292 64218 -71284
rect 68854 -71285 68896 -71272
rect 69202 -71285 69244 -71272
rect 69378 -71274 69440 -71264
rect 69558 -70120 69612 -70110
rect 69558 -71272 69612 -71262
rect 69732 -70118 69794 -70108
rect 69920 -70110 69962 -69842
rect 69732 -71272 69794 -71262
rect 69910 -70120 69964 -70110
rect 70104 -70112 70138 -70094
rect 70278 -70110 70320 -69842
rect 70460 -70104 70494 -70094
rect 69910 -71272 69964 -71262
rect 70094 -70122 70156 -70112
rect 69560 -71275 69602 -71272
rect 69920 -71279 69962 -71272
rect 70094 -71276 70156 -71266
rect 70268 -70120 70322 -70110
rect 70268 -71272 70322 -71262
rect 70452 -70114 70514 -70104
rect 70630 -70110 70672 -69842
rect 70816 -70100 70850 -70094
rect 70804 -70110 70866 -70100
rect 70986 -70104 71028 -69842
rect 71172 -70104 71206 -70094
rect 71344 -70104 71386 -69842
rect 71528 -70104 71562 -70094
rect 70452 -71268 70514 -71258
rect 70620 -70120 70674 -70110
rect 70460 -71270 70494 -71268
rect 70620 -71272 70674 -71262
rect 70804 -71264 70866 -71254
rect 70980 -70114 71034 -70104
rect 70816 -71270 70850 -71264
rect 70980 -71266 71034 -71256
rect 71158 -70114 71220 -70104
rect 70278 -71275 70320 -71272
rect 70630 -71285 70672 -71272
rect 70986 -71285 71028 -71266
rect 71158 -71268 71220 -71258
rect 71336 -70114 71390 -70104
rect 71336 -71266 71390 -71256
rect 71512 -70114 71574 -70104
rect 71700 -70106 71742 -69842
rect 71884 -70104 71918 -70094
rect 71172 -71270 71206 -71268
rect 71344 -71289 71386 -71266
rect 71512 -71268 71574 -71258
rect 71694 -70116 71748 -70106
rect 71694 -71268 71748 -71258
rect 71874 -70114 71936 -70104
rect 72054 -70110 72096 -69842
rect 72240 -70108 72274 -70094
rect 71874 -71268 71936 -71258
rect 72046 -70120 72100 -70110
rect 71528 -71270 71562 -71268
rect 71700 -71285 71742 -71268
rect 71884 -71270 71918 -71268
rect 72046 -71272 72100 -71262
rect 72228 -70118 72290 -70108
rect 72408 -70110 72450 -69842
rect 72596 -70108 72630 -70094
rect 72228 -71272 72290 -71262
rect 72406 -70120 72460 -70110
rect 72406 -71272 72460 -71262
rect 72586 -70118 72648 -70108
rect 72764 -70110 72806 -69842
rect 72952 -70104 72986 -70094
rect 72586 -71272 72648 -71262
rect 72756 -70120 72810 -70110
rect 72756 -71272 72810 -71262
rect 72942 -70114 73004 -70104
rect 73126 -70106 73168 -69842
rect 73308 -70104 73342 -70094
rect 72942 -71268 73004 -71258
rect 73122 -70116 73176 -70106
rect 73122 -71268 73176 -71258
rect 73302 -70114 73364 -70104
rect 73478 -70112 73520 -69842
rect 73664 -70108 73698 -70094
rect 73834 -70106 73876 -69842
rect 74020 -70104 74054 -70094
rect 74190 -70104 74232 -69842
rect 74376 -70102 74410 -70094
rect 73302 -71268 73364 -71258
rect 73472 -70122 73526 -70112
rect 72952 -71270 72986 -71268
rect 72054 -71285 72096 -71272
rect 72408 -71279 72450 -71272
rect 72764 -71289 72806 -71272
rect 73126 -71289 73168 -71268
rect 73308 -71270 73342 -71268
rect 73472 -71274 73526 -71264
rect 73652 -70118 73714 -70108
rect 73652 -71272 73714 -71262
rect 73832 -70116 73886 -70106
rect 73832 -71268 73886 -71258
rect 74008 -70114 74070 -70104
rect 74008 -71268 74070 -71258
rect 74180 -70114 74234 -70104
rect 74180 -71266 74234 -71256
rect 74366 -70112 74428 -70102
rect 74546 -70106 74588 -69842
rect 74732 -70104 74766 -70094
rect 74366 -71266 74428 -71256
rect 74540 -70116 74594 -70106
rect 73478 -71279 73520 -71274
rect 73834 -71289 73876 -71268
rect 74020 -71270 74054 -71268
rect 74190 -71275 74232 -71266
rect 74376 -71270 74410 -71266
rect 74540 -71268 74594 -71258
rect 74724 -70114 74786 -70104
rect 74904 -70106 74946 -69842
rect 75088 -70104 75122 -70094
rect 75258 -70104 75300 -69842
rect 75444 -70102 75478 -70094
rect 74724 -71268 74786 -71258
rect 74896 -70116 74950 -70106
rect 74896 -71268 74950 -71258
rect 75074 -70114 75136 -70104
rect 75074 -71268 75136 -71258
rect 75252 -70114 75306 -70104
rect 75252 -71266 75306 -71256
rect 75432 -70112 75494 -70102
rect 75612 -70106 75654 -69842
rect 75800 -70102 75834 -70094
rect 75972 -70102 76014 -69842
rect 75432 -71266 75494 -71256
rect 75610 -70116 75664 -70106
rect 75258 -71267 75300 -71266
rect 74546 -71285 74588 -71268
rect 74732 -71270 74766 -71268
rect 74904 -71285 74946 -71268
rect 75088 -71270 75122 -71268
rect 75444 -71270 75478 -71266
rect 75610 -71268 75664 -71258
rect 75788 -70112 75850 -70102
rect 75788 -71266 75850 -71256
rect 75966 -70112 76020 -70102
rect 76156 -70104 76190 -70094
rect 75966 -71264 76020 -71254
rect 76146 -70114 76208 -70104
rect 76330 -70106 76372 -69842
rect 76512 -70102 76546 -70094
rect 75612 -71275 75654 -71268
rect 75800 -71270 75834 -71266
rect 75972 -71285 76014 -71264
rect 76146 -71268 76208 -71258
rect 76320 -70116 76374 -70106
rect 76320 -71268 76374 -71258
rect 76496 -70112 76558 -70102
rect 76682 -70106 76724 -69842
rect 76868 -70104 76902 -70094
rect 76496 -71266 76558 -71256
rect 76674 -70116 76728 -70106
rect 76156 -71270 76190 -71268
rect 76330 -71275 76372 -71268
rect 76512 -71270 76546 -71266
rect 76674 -71268 76728 -71258
rect 76860 -70114 76922 -70104
rect 77040 -70106 77082 -69842
rect 76860 -71268 76922 -71258
rect 77036 -70116 77090 -70106
rect 77224 -70108 77258 -70094
rect 77394 -70106 77436 -69842
rect 77580 -70102 77614 -70094
rect 77036 -71268 77090 -71258
rect 77212 -70118 77274 -70108
rect 76682 -71275 76724 -71268
rect 76868 -71270 76902 -71268
rect 77040 -71275 77082 -71268
rect 77212 -71272 77274 -71262
rect 77392 -70116 77446 -70106
rect 77392 -71268 77446 -71258
rect 77568 -70112 77630 -70102
rect 77752 -70110 77794 -69842
rect 77936 -70100 77970 -70094
rect 77926 -70110 77988 -70100
rect 78106 -70106 78148 -69842
rect 78292 -70102 78326 -70094
rect 77568 -71266 77630 -71256
rect 77744 -70120 77798 -70110
rect 77394 -71279 77436 -71268
rect 77580 -71270 77614 -71266
rect 77744 -71272 77798 -71262
rect 77926 -71264 77988 -71254
rect 78104 -70116 78158 -70106
rect 77936 -71270 77970 -71264
rect 78104 -71268 78158 -71258
rect 78282 -70112 78344 -70102
rect 78468 -70106 78510 -69842
rect 78648 -70102 78682 -70094
rect 78282 -71266 78344 -71256
rect 78452 -70116 78510 -70106
rect 78506 -71258 78510 -70116
rect 77752 -71279 77794 -71272
rect 78106 -71275 78148 -71268
rect 78292 -71270 78326 -71266
rect 78452 -71267 78510 -71258
rect 78638 -70112 78700 -70102
rect 78820 -70110 78862 -69842
rect 79004 -70104 79038 -70094
rect 78638 -71266 78700 -71256
rect 78812 -70120 78866 -70110
rect 78452 -71268 78506 -71267
rect 78648 -71270 78682 -71266
rect 78812 -71272 78866 -71262
rect 78996 -70114 79058 -70104
rect 79178 -70106 79220 -69842
rect 78996 -71268 79058 -71258
rect 79170 -70116 79224 -70106
rect 79360 -70108 79394 -70094
rect 79532 -70106 79574 -69842
rect 79170 -71268 79224 -71258
rect 79346 -70118 79408 -70108
rect 79004 -71270 79038 -71268
rect 78820 -71279 78862 -71272
rect 79178 -71275 79220 -71268
rect 79346 -71272 79408 -71262
rect 79522 -70116 79576 -70106
rect 79716 -70108 79750 -70094
rect 79522 -71268 79576 -71258
rect 79704 -70118 79766 -70108
rect 79888 -70110 79930 -69842
rect 80072 -70102 80106 -70094
rect 79704 -71272 79766 -71262
rect 79882 -70120 79936 -70110
rect 79882 -71272 79936 -71262
rect 80058 -70112 80120 -70102
rect 80242 -70106 80284 -69842
rect 80058 -71266 80120 -71256
rect 80236 -70116 80290 -70106
rect 80428 -70108 80462 -70094
rect 80072 -71270 80106 -71266
rect 80236 -71268 80290 -71258
rect 80412 -70118 80474 -70108
rect 80600 -70110 80642 -69842
rect 80784 -70104 80818 -70094
rect 80956 -70104 80998 -69842
rect 79888 -71279 79930 -71272
rect 80242 -71279 80284 -71268
rect 80412 -71272 80474 -71262
rect 80594 -70120 80648 -70110
rect 80594 -71272 80648 -71262
rect 80768 -70114 80830 -70104
rect 80768 -71268 80830 -71258
rect 80948 -70114 81002 -70104
rect 81140 -70108 81174 -70094
rect 81310 -70106 81352 -69842
rect 81496 -70104 81530 -70094
rect 80948 -71266 81002 -71256
rect 81126 -70118 81188 -70108
rect 80784 -71270 80818 -71268
rect 80956 -71275 80998 -71266
rect 81126 -71272 81188 -71262
rect 81306 -70116 81360 -70106
rect 81306 -71268 81360 -71258
rect 81480 -70114 81542 -70104
rect 81666 -70110 81708 -69842
rect 81852 -70108 81886 -70094
rect 81480 -71268 81542 -71258
rect 81660 -70120 81714 -70110
rect 81310 -71279 81352 -71268
rect 81496 -71270 81530 -71268
rect 81660 -71272 81714 -71262
rect 81836 -70118 81898 -70108
rect 82024 -70110 82066 -69842
rect 82208 -70104 82242 -70094
rect 81836 -71272 81898 -71262
rect 82010 -70120 82066 -70110
rect 82064 -71262 82066 -70120
rect 82010 -71272 82066 -71262
rect 82190 -70114 82252 -70104
rect 82382 -70106 82424 -69842
rect 82190 -71268 82252 -71258
rect 82374 -70116 82428 -70106
rect 82564 -70108 82598 -70094
rect 82734 -70106 82776 -69842
rect 82920 -70104 82954 -70094
rect 82374 -71268 82428 -71258
rect 82546 -70118 82608 -70108
rect 82208 -71270 82242 -71268
rect 81666 -71279 81708 -71272
rect 82024 -71275 82066 -71272
rect 82382 -71279 82424 -71268
rect 82546 -71272 82608 -71262
rect 82726 -70116 82780 -70106
rect 82726 -71268 82780 -71258
rect 82906 -70114 82968 -70104
rect 83090 -70106 83132 -69842
rect 83276 -70102 83310 -70094
rect 82906 -71268 82968 -71258
rect 83086 -70116 83140 -70106
rect 83086 -71268 83140 -71258
rect 83264 -70112 83326 -70102
rect 83446 -70112 83488 -69842
rect 83632 -70108 83666 -70094
rect 83264 -71266 83326 -71256
rect 83440 -70122 83494 -70112
rect 82734 -71279 82776 -71268
rect 82920 -71270 82954 -71268
rect 83090 -71289 83132 -71268
rect 83276 -71270 83310 -71266
rect 83440 -71274 83494 -71264
rect 83620 -70118 83682 -70108
rect 83802 -70110 83844 -69842
rect 83988 -70108 84022 -70094
rect 83620 -71272 83682 -71262
rect 83796 -70120 83850 -70110
rect 83796 -71272 83850 -71262
rect 83976 -70118 84038 -70108
rect 84158 -70112 84200 -69842
rect 83976 -71272 84038 -71262
rect 84154 -70122 84208 -70112
rect 64166 -71294 64200 -71292
rect 83446 -71297 83488 -71274
rect 83802 -71285 83844 -71272
rect 84154 -71274 84208 -71264
rect 84158 -71279 84200 -71274
rect 68204 -71328 68302 -71318
rect 60846 -71333 60938 -71330
rect 61202 -71333 61294 -71332
rect 61558 -71333 61650 -71330
rect 61736 -71333 61828 -71330
rect 61916 -71333 62008 -71332
rect 62090 -71333 62182 -71332
rect 62448 -71333 62540 -71332
rect 62810 -71333 62902 -71332
rect 63338 -71333 63430 -71332
rect 63694 -71333 63786 -71332
rect 56330 -71338 59514 -71336
rect 60834 -71338 64295 -71333
rect 68200 -71338 68204 -71328
rect 68374 -71338 68470 -71328
rect 68558 -71338 68654 -71328
rect 68734 -71338 68830 -71328
rect 68912 -71338 69008 -71328
rect 69092 -71338 69188 -71328
rect 69268 -71338 69364 -71328
rect 69444 -71336 69540 -71326
rect 52394 -71340 68200 -71338
rect 52394 -71343 60846 -71340
rect 60938 -71342 61558 -71340
rect 60938 -71343 61202 -71342
rect 61294 -71343 61558 -71342
rect 61650 -71343 61736 -71340
rect 61828 -71342 68200 -71340
rect 61828 -71343 61916 -71342
rect 62008 -71343 62090 -71342
rect 62182 -71343 62448 -71342
rect 62540 -71343 62810 -71342
rect 62902 -71343 63338 -71342
rect 63430 -71343 63694 -71342
rect 63786 -71343 68200 -71342
rect 52394 -71346 60834 -71343
rect 52394 -71478 56330 -71346
rect 59514 -71476 60834 -71346
rect 64295 -71350 68200 -71343
rect 64320 -71406 68200 -71350
rect 59644 -71478 60834 -71476
rect 56330 -71494 59514 -71484
rect 64295 -71478 68200 -71406
rect 60834 -71492 64295 -71482
rect 68302 -71478 68374 -71338
rect 68200 -71492 68204 -71482
rect 68470 -71478 68558 -71338
rect 68374 -71492 68470 -71482
rect 68654 -71478 68734 -71338
rect 68558 -71492 68654 -71482
rect 68830 -71478 68912 -71338
rect 68734 -71492 68830 -71482
rect 69008 -71478 69092 -71338
rect 68912 -71492 69008 -71482
rect 69188 -71478 69268 -71338
rect 69092 -71492 69188 -71482
rect 69364 -71478 69444 -71338
rect 69268 -71492 69364 -71482
rect 69622 -71334 69718 -71324
rect 69540 -71478 69622 -71338
rect 69800 -71336 69896 -71326
rect 69718 -71478 69800 -71338
rect 69444 -71490 69540 -71480
rect 69622 -71488 69718 -71478
rect 69980 -71336 70076 -71326
rect 69896 -71478 69980 -71338
rect 69800 -71490 69896 -71480
rect 70158 -71338 70254 -71328
rect 70338 -71334 70434 -71324
rect 70076 -71478 70158 -71338
rect 69980 -71490 70076 -71480
rect 70254 -71478 70338 -71338
rect 70514 -71338 70610 -71328
rect 70694 -71338 70790 -71328
rect 70874 -71336 70970 -71326
rect 70434 -71478 70514 -71338
rect 70158 -71492 70254 -71482
rect 70338 -71488 70434 -71478
rect 70610 -71478 70694 -71338
rect 70514 -71492 70610 -71482
rect 70790 -71478 70874 -71338
rect 70694 -71492 70790 -71482
rect 71050 -71336 71146 -71326
rect 70970 -71478 71050 -71338
rect 70874 -71490 70970 -71480
rect 71228 -71338 71324 -71328
rect 71404 -71338 71500 -71328
rect 71580 -71336 71676 -71326
rect 71146 -71478 71228 -71338
rect 71050 -71490 71146 -71480
rect 71324 -71478 71404 -71338
rect 71228 -71492 71324 -71482
rect 71500 -71478 71580 -71338
rect 71404 -71492 71500 -71482
rect 71764 -71334 71860 -71324
rect 71676 -71478 71764 -71338
rect 71940 -71338 72036 -71328
rect 72118 -71336 72214 -71326
rect 71860 -71478 71940 -71338
rect 71580 -71490 71676 -71480
rect 71764 -71488 71860 -71478
rect 72036 -71478 72118 -71338
rect 71940 -71492 72036 -71482
rect 72294 -71336 72390 -71326
rect 72214 -71478 72294 -71338
rect 72118 -71490 72214 -71480
rect 72470 -71336 72566 -71326
rect 72390 -71478 72470 -71338
rect 72294 -71490 72390 -71480
rect 72648 -71334 72744 -71324
rect 72566 -71478 72648 -71338
rect 72832 -71336 72928 -71326
rect 72744 -71478 72832 -71338
rect 72470 -71490 72566 -71480
rect 72648 -71488 72744 -71478
rect 73006 -71336 73102 -71326
rect 72928 -71478 73006 -71338
rect 72832 -71490 72928 -71480
rect 73186 -71336 73282 -71326
rect 73102 -71478 73186 -71338
rect 73006 -71490 73102 -71480
rect 73362 -71338 73458 -71328
rect 73542 -71338 73638 -71328
rect 73720 -71338 73816 -71328
rect 73900 -71338 73996 -71328
rect 74074 -71336 74170 -71326
rect 73282 -71478 73362 -71338
rect 73186 -71490 73282 -71480
rect 73458 -71478 73542 -71338
rect 73362 -71492 73458 -71482
rect 73638 -71478 73720 -71338
rect 73542 -71492 73638 -71482
rect 73816 -71478 73900 -71338
rect 73720 -71492 73816 -71482
rect 73996 -71478 74074 -71338
rect 73900 -71492 73996 -71482
rect 74256 -71334 74352 -71324
rect 74170 -71478 74256 -71338
rect 74434 -71336 74530 -71326
rect 74352 -71478 74434 -71338
rect 74074 -71490 74170 -71480
rect 74256 -71488 74352 -71478
rect 74614 -71334 74710 -71324
rect 74530 -71478 74614 -71338
rect 74792 -71332 74888 -71322
rect 74710 -71476 74792 -71338
rect 74968 -71334 75064 -71324
rect 74888 -71476 74968 -71338
rect 74710 -71478 74968 -71476
rect 75146 -71336 75242 -71326
rect 75064 -71478 75146 -71338
rect 74434 -71490 74530 -71480
rect 74614 -71488 74710 -71478
rect 74792 -71486 74888 -71478
rect 74968 -71488 75064 -71478
rect 75326 -71334 75422 -71324
rect 75242 -71478 75326 -71338
rect 75502 -71338 75598 -71328
rect 75680 -71334 75776 -71324
rect 75422 -71478 75502 -71338
rect 75146 -71490 75242 -71480
rect 75326 -71488 75422 -71478
rect 75598 -71478 75680 -71338
rect 75856 -71334 75952 -71324
rect 75776 -71478 75856 -71338
rect 76034 -71334 76130 -71324
rect 75952 -71478 76034 -71338
rect 76214 -71334 76310 -71324
rect 76130 -71478 76214 -71338
rect 76392 -71336 76488 -71326
rect 76310 -71478 76392 -71338
rect 75502 -71492 75598 -71482
rect 75680 -71488 75776 -71478
rect 75856 -71488 75952 -71478
rect 76034 -71488 76130 -71478
rect 76214 -71488 76310 -71478
rect 76572 -71334 76668 -71324
rect 76488 -71478 76572 -71338
rect 76746 -71336 76842 -71326
rect 76668 -71478 76746 -71338
rect 76392 -71490 76488 -71480
rect 76572 -71488 76668 -71478
rect 76922 -71336 77018 -71326
rect 76842 -71478 76922 -71338
rect 76746 -71490 76842 -71480
rect 77102 -71336 77198 -71326
rect 77018 -71478 77102 -71338
rect 76922 -71490 77018 -71480
rect 77282 -71336 77378 -71326
rect 77198 -71478 77282 -71338
rect 77102 -71490 77198 -71480
rect 77458 -71338 77554 -71328
rect 77636 -71336 77732 -71326
rect 77378 -71478 77458 -71338
rect 77282 -71490 77378 -71480
rect 77554 -71478 77636 -71338
rect 77458 -71492 77554 -71482
rect 77814 -71336 77910 -71326
rect 77732 -71478 77814 -71338
rect 77636 -71490 77732 -71480
rect 77990 -71334 78086 -71324
rect 77910 -71478 77990 -71338
rect 78168 -71334 78264 -71324
rect 78086 -71478 78168 -71338
rect 78348 -71334 78444 -71324
rect 78264 -71478 78348 -71338
rect 78526 -71334 78622 -71324
rect 78444 -71478 78526 -71338
rect 78704 -71334 78800 -71324
rect 78622 -71478 78704 -71338
rect 78882 -71334 78978 -71324
rect 78800 -71478 78882 -71338
rect 79062 -71334 79158 -71324
rect 78978 -71478 79062 -71338
rect 79236 -71336 79332 -71326
rect 79158 -71478 79236 -71338
rect 77814 -71490 77910 -71480
rect 77990 -71488 78086 -71478
rect 78168 -71488 78264 -71478
rect 78348 -71488 78444 -71478
rect 78526 -71488 78622 -71478
rect 78704 -71488 78800 -71478
rect 78882 -71488 78978 -71478
rect 79062 -71488 79158 -71478
rect 79412 -71338 79508 -71328
rect 79592 -71336 79688 -71326
rect 79332 -71478 79412 -71338
rect 79236 -71490 79332 -71480
rect 79508 -71478 79592 -71338
rect 79412 -71492 79508 -71482
rect 79770 -71336 79866 -71326
rect 79688 -71478 79770 -71338
rect 79592 -71490 79688 -71480
rect 79948 -71336 80044 -71326
rect 79866 -71478 79948 -71338
rect 79770 -71490 79866 -71480
rect 80126 -71336 80222 -71326
rect 80044 -71478 80126 -71338
rect 79948 -71490 80044 -71480
rect 80304 -71336 80400 -71326
rect 80222 -71478 80304 -71338
rect 80126 -71490 80222 -71480
rect 80484 -71336 80580 -71326
rect 80400 -71478 80484 -71338
rect 80304 -71490 80400 -71480
rect 80662 -71336 80758 -71326
rect 80580 -71478 80662 -71338
rect 80484 -71490 80580 -71480
rect 80840 -71334 80936 -71324
rect 80758 -71478 80840 -71338
rect 81016 -71334 81112 -71324
rect 80936 -71478 81016 -71338
rect 81198 -71334 81294 -71324
rect 81112 -71478 81198 -71338
rect 81372 -71334 81468 -71324
rect 81294 -71478 81372 -71338
rect 81554 -71334 81650 -71324
rect 81468 -71478 81554 -71338
rect 81732 -71336 81828 -71326
rect 81650 -71478 81732 -71338
rect 80662 -71490 80758 -71480
rect 80840 -71488 80936 -71478
rect 81016 -71488 81112 -71478
rect 81198 -71488 81294 -71478
rect 81372 -71488 81468 -71478
rect 81554 -71488 81650 -71478
rect 81908 -71336 82004 -71326
rect 81828 -71478 81908 -71338
rect 81732 -71490 81828 -71480
rect 82086 -71334 82182 -71324
rect 82004 -71478 82086 -71338
rect 82264 -71334 82360 -71324
rect 82182 -71478 82264 -71338
rect 82444 -71336 82540 -71326
rect 82360 -71478 82444 -71338
rect 81908 -71490 82004 -71480
rect 82086 -71488 82182 -71478
rect 82264 -71488 82360 -71478
rect 82622 -71336 82718 -71326
rect 82540 -71478 82622 -71338
rect 82444 -71490 82540 -71480
rect 82798 -71336 82894 -71326
rect 82718 -71478 82798 -71338
rect 82622 -71490 82718 -71480
rect 82980 -71336 83076 -71326
rect 82894 -71478 82980 -71338
rect 82798 -71490 82894 -71480
rect 83158 -71336 83254 -71326
rect 83076 -71478 83158 -71338
rect 82980 -71490 83076 -71480
rect 83334 -71334 83430 -71324
rect 83254 -71478 83334 -71338
rect 83512 -71334 83608 -71324
rect 83430 -71478 83512 -71338
rect 83688 -71334 83784 -71324
rect 83608 -71478 83688 -71338
rect 83868 -71336 83964 -71326
rect 83784 -71478 83868 -71338
rect 83158 -71490 83254 -71480
rect 83334 -71488 83430 -71478
rect 83512 -71488 83608 -71478
rect 83688 -71488 83784 -71478
rect 84046 -71336 84142 -71326
rect 83964 -71478 84046 -71338
rect 83868 -71490 83964 -71480
rect 84142 -71478 84258 -71338
rect 84046 -71490 84142 -71480
rect 68204 -71502 68302 -71492
rect 68136 -71552 68178 -71536
rect 68322 -71552 68356 -71536
rect 68488 -71544 68530 -71536
rect 68664 -71540 68726 -71530
rect 68132 -71562 68190 -71552
rect 56242 -73154 66630 -72608
rect 68132 -72716 68190 -72706
rect 68314 -71562 68376 -71552
rect 68314 -72716 68376 -72706
rect 68488 -71554 68552 -71544
rect 68488 -72698 68494 -71554
rect 68852 -71544 68894 -71536
rect 69018 -71542 69080 -71532
rect 68664 -72694 68668 -72684
rect 68488 -72708 68552 -72698
rect 68668 -72708 68726 -72698
rect 68848 -71554 68906 -71544
rect 69080 -71554 69086 -71544
rect 69018 -72662 69028 -72652
rect 68848 -72708 68906 -72698
rect 69028 -72708 69086 -72698
rect 69200 -71546 69242 -71536
rect 69378 -71540 69440 -71530
rect 70086 -71536 70148 -71526
rect 69200 -71556 69260 -71546
rect 69200 -72700 69202 -71556
rect 69558 -71544 69600 -71536
rect 69746 -71538 69780 -71536
rect 69378 -72694 69382 -72684
rect 68136 -72930 68178 -72716
rect 68488 -72930 68530 -72708
rect 68678 -72712 68712 -72708
rect 68852 -72930 68894 -72708
rect 69034 -72712 69068 -72708
rect 69200 -72710 69260 -72700
rect 69200 -72930 69242 -72710
rect 69382 -72712 69440 -72702
rect 69556 -71554 69614 -71544
rect 69724 -71548 69786 -71538
rect 69918 -71550 69960 -71536
rect 69786 -71562 69798 -71552
rect 69724 -72668 69740 -72658
rect 69556 -72708 69614 -72698
rect 69558 -72930 69600 -72708
rect 69740 -72716 69798 -72706
rect 69910 -71560 69968 -71550
rect 70148 -71560 70150 -71550
rect 70276 -71552 70318 -71536
rect 70450 -71542 70512 -71532
rect 70086 -72656 70092 -72646
rect 69910 -72714 69968 -72704
rect 70092 -72714 70150 -72704
rect 70266 -71562 70324 -71552
rect 69918 -72930 69960 -72714
rect 70266 -72716 70324 -72706
rect 70444 -71560 70450 -71550
rect 70628 -71548 70670 -71536
rect 70790 -71546 70852 -71536
rect 70984 -71546 71026 -71537
rect 71170 -71544 71204 -71536
rect 70502 -72662 70512 -72652
rect 70624 -71558 70682 -71548
rect 70444 -72714 70502 -72704
rect 70852 -71560 70858 -71550
rect 70790 -72666 70800 -72656
rect 70624 -72712 70682 -72702
rect 70276 -72930 70318 -72716
rect 70628 -72930 70670 -72712
rect 70800 -72714 70858 -72704
rect 70982 -71556 71040 -71546
rect 71148 -71548 71210 -71544
rect 71148 -71554 71214 -71548
rect 71342 -71550 71384 -71537
rect 71504 -71546 71566 -71536
rect 71210 -71558 71214 -71554
rect 71148 -72674 71156 -72664
rect 70982 -72710 71040 -72700
rect 70984 -72930 71026 -72710
rect 71156 -72712 71214 -72702
rect 71336 -71560 71394 -71550
rect 71566 -71558 71574 -71548
rect 71698 -71550 71740 -71536
rect 71858 -71542 71920 -71532
rect 71504 -72666 71516 -72656
rect 71336 -72714 71394 -72704
rect 71516 -72712 71574 -72702
rect 71692 -71560 71750 -71550
rect 72052 -71548 72094 -71536
rect 72216 -71546 72278 -71536
rect 71920 -71558 71928 -71548
rect 71858 -72662 71870 -72652
rect 71692 -72714 71750 -72704
rect 71870 -72712 71928 -72702
rect 72048 -71558 72106 -71548
rect 72278 -71558 72288 -71548
rect 72406 -71552 72448 -71539
rect 72570 -71544 72632 -71534
rect 72216 -72666 72230 -72656
rect 72048 -72712 72106 -72702
rect 72230 -72712 72288 -72702
rect 72404 -71562 72462 -71552
rect 72762 -71550 72804 -71537
rect 72946 -71542 73008 -71532
rect 73988 -71536 74050 -71532
rect 75764 -71536 75826 -71534
rect 72632 -71560 72644 -71550
rect 72570 -72664 72586 -72654
rect 71342 -72930 71384 -72714
rect 71698 -72930 71740 -72714
rect 72052 -72930 72094 -72712
rect 72404 -72716 72462 -72706
rect 72586 -72714 72644 -72704
rect 72754 -71560 72812 -71550
rect 72754 -72714 72812 -72704
rect 72938 -71558 72946 -71548
rect 73124 -71548 73166 -71537
rect 73306 -71548 73340 -71536
rect 73476 -71546 73518 -71536
rect 73662 -71540 73696 -71536
rect 72996 -72662 73008 -72652
rect 73118 -71558 73176 -71548
rect 72938 -72712 72996 -72702
rect 73286 -71552 73348 -71548
rect 73286 -71558 73350 -71552
rect 73348 -71562 73350 -71558
rect 73286 -72678 73292 -72668
rect 73118 -72712 73176 -72702
rect 72406 -72930 72448 -72716
rect 72762 -72930 72804 -72714
rect 73124 -72930 73166 -72712
rect 73292 -72716 73350 -72706
rect 73466 -71556 73524 -71546
rect 73642 -71550 73704 -71540
rect 73832 -71544 73874 -71539
rect 73988 -71542 74052 -71536
rect 73704 -71560 73712 -71550
rect 73642 -72670 73654 -72660
rect 73466 -72710 73524 -72700
rect 73476 -72930 73518 -72710
rect 73654 -72714 73712 -72704
rect 73830 -71554 73888 -71544
rect 74050 -71544 74052 -71542
rect 74050 -71554 74068 -71544
rect 73988 -72662 74010 -72652
rect 73830 -72708 73888 -72698
rect 74010 -72708 74068 -72698
rect 74188 -71546 74230 -71536
rect 74374 -71542 74408 -71536
rect 74544 -71542 74586 -71539
rect 74188 -71556 74246 -71546
rect 74364 -71550 74422 -71542
rect 74352 -71552 74422 -71550
rect 74352 -71560 74364 -71552
rect 74352 -72680 74364 -72670
rect 73832 -72930 73874 -72708
rect 74018 -72712 74052 -72708
rect 74188 -72710 74246 -72700
rect 74364 -72706 74422 -72696
rect 74544 -71552 74602 -71542
rect 74730 -71544 74764 -71536
rect 74902 -71544 74944 -71536
rect 74720 -71546 74778 -71544
rect 74714 -71554 74778 -71546
rect 74714 -71556 74720 -71554
rect 74714 -72676 74720 -72666
rect 74544 -72706 74602 -72696
rect 74188 -72930 74230 -72710
rect 74374 -72712 74408 -72706
rect 74544 -72930 74586 -72706
rect 74720 -72708 74778 -72698
rect 74898 -71554 74956 -71544
rect 75086 -71554 75120 -71536
rect 75256 -71552 75298 -71536
rect 75442 -71548 75476 -71536
rect 75432 -71550 75490 -71548
rect 75078 -71562 75136 -71554
rect 75068 -71564 75136 -71562
rect 75068 -71572 75078 -71564
rect 75068 -72692 75078 -72682
rect 74898 -72708 74956 -72698
rect 74730 -72712 74764 -72708
rect 74902 -72930 74944 -72708
rect 75078 -72718 75136 -72708
rect 75246 -71562 75304 -71552
rect 75426 -71558 75490 -71550
rect 75426 -71560 75432 -71558
rect 75610 -71562 75652 -71539
rect 75764 -71544 75832 -71536
rect 75426 -72680 75432 -72670
rect 75246 -72716 75304 -72706
rect 75432 -72712 75490 -72702
rect 75608 -71572 75666 -71562
rect 75826 -71554 75832 -71544
rect 75970 -71554 76012 -71537
rect 76130 -71542 76192 -71532
rect 76478 -71536 76540 -71532
rect 76328 -71542 76370 -71537
rect 76478 -71542 76544 -71536
rect 75826 -71564 75844 -71554
rect 75764 -72664 75786 -72654
rect 75256 -72930 75298 -72716
rect 75608 -72726 75666 -72716
rect 75786 -72718 75844 -72708
rect 75964 -71564 76022 -71554
rect 76192 -71556 76204 -71546
rect 76130 -72662 76146 -72652
rect 75964 -72718 76022 -72708
rect 76146 -72710 76204 -72700
rect 76326 -71552 76384 -71542
rect 76540 -71546 76544 -71542
rect 76540 -71556 76558 -71546
rect 76680 -71552 76722 -71537
rect 76854 -71546 76916 -71536
rect 76478 -72662 76500 -72652
rect 76326 -72706 76384 -72696
rect 76154 -72712 76188 -72710
rect 75610 -72930 75652 -72726
rect 75970 -72930 76012 -72718
rect 76328 -72930 76370 -72706
rect 76500 -72710 76558 -72700
rect 76674 -71562 76732 -71552
rect 76510 -72712 76544 -72710
rect 76674 -72716 76732 -72706
rect 77038 -71550 77080 -71536
rect 77222 -71540 77256 -71536
rect 77196 -71550 77258 -71540
rect 76912 -72666 76916 -72656
rect 77034 -71560 77092 -71550
rect 76854 -72716 76912 -72706
rect 77258 -71562 77270 -71552
rect 77392 -71554 77434 -71536
rect 77578 -71552 77612 -71536
rect 77750 -71548 77792 -71536
rect 77908 -71538 77970 -71528
rect 77196 -72670 77212 -72660
rect 77034 -72714 77092 -72704
rect 76680 -72930 76722 -72716
rect 77038 -72930 77080 -72714
rect 77212 -72716 77270 -72706
rect 77386 -71564 77444 -71554
rect 77548 -71562 77624 -71552
rect 77548 -72682 77566 -72672
rect 77386 -72718 77444 -72708
rect 77566 -72716 77624 -72706
rect 77744 -71558 77802 -71548
rect 78104 -71552 78146 -71536
rect 78274 -71540 78336 -71530
rect 77970 -71564 77982 -71554
rect 77908 -72658 77924 -72648
rect 77744 -72712 77802 -72702
rect 77392 -72930 77434 -72718
rect 77750 -72930 77792 -72712
rect 77924 -72718 77982 -72708
rect 78104 -71562 78162 -71552
rect 78466 -71560 78508 -71539
rect 78646 -71552 78680 -71536
rect 78818 -71552 78860 -71536
rect 79002 -71552 79036 -71536
rect 78624 -71558 78686 -71552
rect 78274 -72660 78276 -72650
rect 78104 -72716 78162 -72706
rect 78334 -72660 78336 -72650
rect 78458 -71570 78516 -71560
rect 78104 -72930 78146 -72716
rect 78276 -72722 78334 -72712
rect 78624 -71562 78694 -71558
rect 78686 -71568 78694 -71562
rect 78624 -72682 78636 -72672
rect 78458 -72724 78516 -72714
rect 78636 -72722 78694 -72712
rect 78810 -71562 78868 -71552
rect 78810 -72716 78868 -72706
rect 78990 -71562 79052 -71552
rect 79176 -71554 79218 -71536
rect 79338 -71542 79400 -71532
rect 79048 -72682 79052 -72672
rect 79170 -71564 79228 -71554
rect 78466 -72930 78508 -72724
rect 78818 -72930 78860 -72716
rect 78990 -72722 79048 -72712
rect 79530 -71552 79572 -71536
rect 79714 -71540 79748 -71536
rect 79692 -71550 79754 -71540
rect 79886 -71550 79928 -71537
rect 80070 -71546 80104 -71536
rect 80048 -71550 80110 -71546
rect 80240 -71550 80282 -71537
rect 80426 -71548 80460 -71536
rect 80598 -71546 80640 -71539
rect 80782 -71542 80816 -71536
rect 80416 -71550 80474 -71548
rect 79400 -71566 79402 -71556
rect 79338 -72662 79344 -72652
rect 79170 -72718 79228 -72708
rect 79176 -72930 79218 -72718
rect 79344 -72720 79402 -72710
rect 79526 -71562 79584 -71552
rect 79754 -71562 79758 -71552
rect 79692 -72670 79700 -72660
rect 79526 -72716 79584 -72706
rect 79700 -72716 79758 -72706
rect 79882 -71560 79940 -71550
rect 80048 -71556 80116 -71550
rect 80110 -71560 80116 -71556
rect 80048 -72676 80058 -72666
rect 79882 -72714 79940 -72704
rect 80058 -72714 80116 -72704
rect 80232 -71560 80290 -71550
rect 80398 -71558 80474 -71550
rect 80398 -71560 80416 -71558
rect 80398 -72680 80416 -72670
rect 80232 -72714 80290 -72704
rect 80416 -72712 80474 -72702
rect 80590 -71556 80648 -71546
rect 80760 -71552 80822 -71542
rect 80954 -71548 80996 -71539
rect 80822 -71562 80830 -71552
rect 80760 -72672 80772 -72662
rect 80590 -72710 80648 -72700
rect 79530 -72930 79572 -72716
rect 79886 -72930 79928 -72714
rect 80240 -72930 80282 -72714
rect 80598 -72930 80640 -72710
rect 80772 -72716 80830 -72706
rect 80946 -71558 81004 -71548
rect 81138 -71550 81172 -71536
rect 81308 -71546 81350 -71537
rect 81494 -71540 81528 -71536
rect 81124 -71552 81182 -71550
rect 81120 -71560 81182 -71552
rect 81120 -71562 81124 -71560
rect 81120 -72682 81124 -72672
rect 80946 -72712 81004 -72702
rect 80954 -72930 80996 -72712
rect 81124 -72714 81182 -72704
rect 81298 -71556 81356 -71546
rect 81478 -71550 81540 -71540
rect 81664 -71546 81706 -71536
rect 81850 -71542 81884 -71536
rect 81848 -71546 81910 -71542
rect 81478 -72670 81482 -72660
rect 81298 -72710 81356 -72700
rect 81482 -72710 81540 -72700
rect 81658 -71556 81716 -71546
rect 81658 -72710 81716 -72700
rect 81836 -71552 81910 -71546
rect 82022 -71548 82064 -71537
rect 81836 -71556 81848 -71552
rect 81894 -72672 81910 -72662
rect 82018 -71558 82076 -71548
rect 82206 -71550 82240 -71536
rect 81836 -72710 81894 -72700
rect 82186 -71560 82254 -71550
rect 82380 -71552 82422 -71536
rect 82562 -71548 82596 -71536
rect 82186 -72680 82196 -72670
rect 81308 -72930 81350 -72710
rect 81494 -72712 81528 -72710
rect 81664 -72930 81706 -72710
rect 81850 -72712 81884 -72710
rect 82018 -72712 82076 -72702
rect 82022 -72930 82064 -72712
rect 82196 -72714 82254 -72704
rect 82370 -71562 82428 -71552
rect 82556 -71556 82614 -71548
rect 82732 -71550 82774 -71536
rect 82918 -71544 82952 -71536
rect 83088 -71544 83130 -71536
rect 83274 -71542 83308 -71536
rect 82542 -71558 82614 -71556
rect 82542 -71566 82556 -71558
rect 82542 -72686 82556 -72676
rect 82370 -72716 82428 -72706
rect 82556 -72712 82614 -72702
rect 82724 -71560 82782 -71550
rect 82724 -72714 82782 -72704
rect 82908 -71554 82966 -71544
rect 83080 -71554 83138 -71544
rect 82966 -71574 82972 -71564
rect 82966 -72694 82972 -72684
rect 82908 -72708 82966 -72698
rect 83258 -71552 83320 -71542
rect 83258 -72672 83262 -72662
rect 83080 -72708 83138 -72698
rect 83262 -72708 83320 -72698
rect 83444 -71550 83486 -71536
rect 83444 -71560 83502 -71550
rect 83630 -71552 83664 -71536
rect 83800 -71552 83842 -71536
rect 83986 -71540 84020 -71536
rect 83962 -71546 84024 -71540
rect 83962 -71550 84036 -71546
rect 83622 -71562 83680 -71552
rect 83612 -71574 83622 -71564
rect 83612 -72694 83622 -72684
rect 82918 -72712 82952 -72708
rect 82380 -72930 82422 -72716
rect 82732 -72930 82774 -72714
rect 83088 -72930 83130 -72708
rect 83274 -72712 83308 -72708
rect 83444 -72714 83502 -72704
rect 83444 -72930 83486 -72714
rect 83622 -72716 83680 -72706
rect 83796 -71562 83854 -71552
rect 84024 -71556 84036 -71550
rect 84156 -71556 84198 -71536
rect 83962 -72670 83978 -72660
rect 83796 -72716 83854 -72706
rect 83978 -72710 84036 -72700
rect 84148 -71566 84206 -71556
rect 83986 -72712 84020 -72710
rect 83800 -72930 83842 -72716
rect 84148 -72720 84206 -72710
rect 84156 -72930 84198 -72720
rect 84320 -72930 86894 -69842
rect 56300 -73388 56354 -73154
rect 56502 -73386 56536 -73378
rect 56300 -73398 56368 -73388
rect 56490 -73392 56544 -73386
rect 56300 -74539 56314 -73398
rect 56314 -74554 56368 -74544
rect 56488 -73396 56544 -73392
rect 56488 -73402 56490 -73396
rect 56488 -74542 56490 -74540
rect 56488 -74550 56544 -74542
rect 56490 -74552 56544 -74550
rect 56654 -73390 56708 -73154
rect 56858 -73386 56892 -73376
rect 56654 -73400 56722 -73390
rect 56654 -74546 56668 -73400
rect 56502 -74554 56536 -74552
rect 56654 -74556 56722 -74546
rect 56852 -73396 56908 -73386
rect 56906 -74542 56908 -74534
rect 56852 -74544 56908 -74542
rect 57010 -73394 57064 -73154
rect 57010 -73404 57080 -73394
rect 57214 -73398 57248 -73376
rect 57368 -73394 57422 -73154
rect 57570 -73390 57604 -73376
rect 57718 -73390 57772 -73154
rect 57558 -73392 57612 -73390
rect 56852 -74552 56906 -74544
rect 57010 -74550 57026 -73404
rect 57010 -74555 57080 -74550
rect 56654 -74559 56708 -74556
rect 57026 -74560 57080 -74555
rect 57196 -73408 57256 -73398
rect 57196 -74554 57202 -74546
rect 57196 -74556 57256 -74554
rect 57368 -73404 57436 -73394
rect 57368 -74550 57382 -73404
rect 57556 -73400 57612 -73392
rect 57556 -73402 57558 -73400
rect 57556 -74546 57558 -74540
rect 57556 -74550 57612 -74546
rect 57368 -74555 57436 -74550
rect 57202 -74564 57256 -74556
rect 57382 -74560 57436 -74555
rect 57558 -74556 57612 -74550
rect 57718 -73400 57794 -73390
rect 57924 -73394 57958 -73378
rect 58082 -73394 58136 -73154
rect 57718 -74546 57740 -73400
rect 57718 -74555 57794 -74546
rect 57740 -74556 57794 -74555
rect 57916 -73398 57970 -73394
rect 57916 -73404 57972 -73398
rect 57970 -73408 57972 -73404
rect 57970 -74550 57972 -74546
rect 57916 -74556 57972 -74550
rect 58082 -73404 58148 -73394
rect 58282 -73398 58316 -73376
rect 58432 -73394 58486 -73154
rect 58638 -73390 58672 -73376
rect 58276 -73400 58330 -73398
rect 58082 -74550 58094 -73404
rect 58082 -74555 58148 -74550
rect 57916 -74560 57970 -74556
rect 58094 -74560 58148 -74555
rect 58274 -73408 58330 -73400
rect 58274 -73410 58276 -73408
rect 58274 -74554 58276 -74548
rect 58274 -74558 58330 -74554
rect 58276 -74564 58330 -74558
rect 58432 -73404 58504 -73394
rect 58432 -74550 58450 -73404
rect 58628 -73400 58684 -73390
rect 58628 -74548 58630 -74538
rect 58432 -74559 58504 -74550
rect 58630 -74558 58684 -74548
rect 58790 -73392 58844 -73154
rect 58994 -73390 59028 -73378
rect 59146 -73390 59200 -73154
rect 59350 -73390 59384 -73376
rect 59496 -73386 59550 -73154
rect 58790 -73402 58860 -73392
rect 58986 -73394 59040 -73390
rect 58790 -74548 58806 -73402
rect 58790 -74555 58860 -74548
rect 58980 -73400 59040 -73394
rect 58980 -73404 58986 -73400
rect 58980 -74546 58986 -74542
rect 58980 -74552 59040 -74546
rect 58806 -74558 58860 -74555
rect 58986 -74556 59040 -74552
rect 59146 -73400 59220 -73390
rect 59146 -74546 59166 -73400
rect 59146 -74556 59220 -74546
rect 59342 -73400 59398 -73390
rect 59342 -74546 59344 -74538
rect 59342 -74548 59398 -74546
rect 59344 -74556 59398 -74548
rect 59496 -73396 59576 -73386
rect 59706 -73390 59740 -73376
rect 59698 -73394 59752 -73390
rect 59496 -74542 59522 -73396
rect 59496 -74552 59576 -74542
rect 59694 -73400 59752 -73394
rect 59694 -73404 59698 -73400
rect 59694 -74546 59698 -74542
rect 59694 -74552 59752 -74546
rect 59496 -74555 59550 -74552
rect 59698 -74556 59752 -74552
rect 59862 -73394 59916 -73154
rect 60062 -73394 60096 -73378
rect 60208 -73394 60262 -73154
rect 59862 -73404 59930 -73394
rect 60054 -73402 60108 -73394
rect 59862 -74550 59876 -73404
rect 59862 -74555 59930 -74550
rect 59146 -74559 59200 -74556
rect 58450 -74560 58504 -74559
rect 59876 -74560 59930 -74555
rect 60052 -73404 60108 -73402
rect 60052 -73412 60054 -73404
rect 60052 -74560 60108 -74550
rect 60208 -73404 60282 -73394
rect 60418 -73398 60452 -73380
rect 60568 -73398 60622 -73154
rect 60774 -73390 60808 -73380
rect 60768 -73396 60822 -73390
rect 60406 -73400 60460 -73398
rect 60208 -74550 60228 -73404
rect 60208 -74559 60282 -74550
rect 60402 -73408 60460 -73400
rect 60402 -73410 60406 -73408
rect 60402 -74554 60406 -74548
rect 60402 -74558 60460 -74554
rect 60228 -74560 60282 -74559
rect 60406 -74564 60460 -74558
rect 60568 -73408 60642 -73398
rect 60568 -74554 60588 -73408
rect 60764 -73400 60822 -73396
rect 60764 -73406 60768 -73400
rect 60764 -74546 60768 -74544
rect 60764 -74554 60822 -74546
rect 60568 -74564 60642 -74554
rect 60768 -74556 60822 -74554
rect 60926 -73394 60980 -73154
rect 61130 -73394 61164 -73380
rect 60926 -73404 60998 -73394
rect 61122 -73400 61176 -73394
rect 60926 -74550 60944 -73404
rect 60926 -74559 60998 -74550
rect 61118 -73404 61176 -73400
rect 61118 -73410 61122 -73404
rect 61118 -74550 61122 -74548
rect 61118 -74558 61176 -74550
rect 61280 -73398 61334 -73154
rect 61486 -73392 61520 -73380
rect 61636 -73390 61690 -73154
rect 61478 -73394 61532 -73392
rect 61280 -73408 61352 -73398
rect 61280 -74554 61298 -73408
rect 61476 -73402 61532 -73394
rect 61476 -73404 61478 -73402
rect 61476 -74548 61478 -74542
rect 61476 -74552 61532 -74548
rect 61280 -74555 61352 -74554
rect 60944 -74560 60998 -74559
rect 61122 -74560 61176 -74558
rect 61298 -74564 61352 -74555
rect 61478 -74558 61532 -74552
rect 61636 -73400 61710 -73390
rect 61842 -73394 61876 -73382
rect 61994 -73394 62048 -73154
rect 62198 -73394 62232 -73384
rect 62352 -73394 62406 -73154
rect 62554 -73392 62588 -73380
rect 62708 -73388 62762 -73154
rect 61828 -73400 61882 -73394
rect 61636 -74546 61656 -73400
rect 61636 -74555 61710 -74546
rect 61656 -74556 61710 -74555
rect 61826 -73404 61882 -73400
rect 61826 -73410 61828 -73404
rect 61826 -74550 61828 -74548
rect 61826 -74558 61882 -74550
rect 61828 -74560 61882 -74558
rect 61994 -73404 62062 -73394
rect 61994 -74550 62008 -73404
rect 61994 -74559 62062 -74550
rect 62008 -74560 62062 -74559
rect 62188 -73404 62242 -73394
rect 62352 -73404 62422 -73394
rect 62546 -73400 62600 -73392
rect 62242 -73414 62244 -73404
rect 62188 -74562 62244 -74552
rect 62352 -74550 62368 -73404
rect 62352 -74555 62422 -74550
rect 62368 -74560 62422 -74555
rect 62544 -73402 62600 -73400
rect 62544 -73410 62546 -73402
rect 62544 -74558 62600 -74548
rect 62708 -73398 62774 -73388
rect 62910 -73394 62944 -73378
rect 63058 -73392 63112 -73154
rect 63266 -73388 63300 -73378
rect 62708 -74544 62720 -73398
rect 62898 -73404 62952 -73394
rect 62708 -74554 62774 -74544
rect 62894 -73414 62898 -73404
rect 62950 -74552 62952 -74550
rect 62708 -74559 62762 -74554
rect 62894 -74560 62952 -74552
rect 63058 -73402 63134 -73392
rect 63256 -73398 63310 -73388
rect 63058 -74548 63080 -73402
rect 63058 -74558 63134 -74548
rect 63254 -73412 63256 -73402
rect 62894 -74562 62950 -74560
rect 60568 -74571 60622 -74564
rect 63058 -74571 63112 -74558
rect 63254 -74560 63310 -74550
rect 63416 -73392 63470 -73154
rect 63622 -73390 63656 -73378
rect 63774 -73390 63828 -73154
rect 63978 -73388 64012 -73378
rect 64126 -73386 64180 -73154
rect 63416 -73402 63486 -73392
rect 63416 -74548 63432 -73402
rect 63416 -74558 63486 -74548
rect 63612 -73400 63666 -73390
rect 63774 -73400 63844 -73390
rect 63968 -73398 64022 -73388
rect 63666 -73414 63670 -73404
rect 63612 -74552 63614 -74546
rect 63612 -74556 63670 -74552
rect 63774 -74546 63790 -73400
rect 63774 -74555 63844 -74546
rect 63790 -74556 63844 -74555
rect 63966 -73408 63968 -73398
rect 64126 -73396 64200 -73386
rect 64334 -73390 64368 -73380
rect 64126 -74539 64146 -73396
rect 63966 -74556 64022 -74546
rect 64322 -73398 64376 -73390
rect 64146 -74552 64200 -74542
rect 64320 -73400 64376 -73398
rect 64320 -73408 64322 -73400
rect 64320 -74556 64376 -74546
rect 63416 -74559 63470 -74558
rect 63614 -74562 63670 -74556
rect 56364 -74628 56470 -74626
rect 57086 -74628 57192 -74626
rect 57262 -74628 57368 -74626
rect 59390 -74628 59496 -74626
rect 59568 -74628 59674 -74622
rect 62240 -74628 62346 -74622
rect 63848 -74628 63954 -74626
rect 64200 -74628 64306 -74626
rect 54812 -74632 64372 -74628
rect 54812 -74636 59568 -74632
rect 54812 -74792 56364 -74636
rect 56470 -74638 57086 -74636
rect 56470 -74642 56728 -74638
rect 56470 -74792 56546 -74642
rect 54812 -74796 56546 -74792
rect 54815 -76432 54962 -74796
rect 56364 -74802 56470 -74796
rect 56652 -74794 56728 -74642
rect 56834 -74794 56908 -74638
rect 57014 -74792 57086 -74638
rect 57192 -74792 57262 -74636
rect 57368 -74638 59390 -74636
rect 57368 -74792 57446 -74638
rect 57014 -74794 57446 -74792
rect 57552 -74794 57620 -74638
rect 57726 -74794 57794 -74638
rect 57900 -74642 58150 -74638
rect 57900 -74794 57976 -74642
rect 56652 -74796 57976 -74794
rect 56546 -74808 56652 -74798
rect 56728 -74804 56834 -74796
rect 56908 -74804 57014 -74796
rect 57086 -74802 57192 -74796
rect 57262 -74802 57368 -74796
rect 57446 -74804 57552 -74796
rect 57620 -74804 57726 -74796
rect 57794 -74804 57900 -74796
rect 58082 -74794 58150 -74642
rect 58256 -74794 58328 -74638
rect 58434 -74794 58508 -74638
rect 58614 -74794 58678 -74638
rect 58784 -74794 58858 -74638
rect 58964 -74794 59042 -74638
rect 59148 -74794 59216 -74638
rect 59322 -74792 59390 -74638
rect 59496 -74788 59568 -74636
rect 59674 -74638 62240 -74632
rect 59674 -74642 59926 -74638
rect 59674 -74788 59750 -74642
rect 59496 -74792 59750 -74788
rect 59322 -74794 59750 -74792
rect 58082 -74796 59750 -74794
rect 57976 -74808 58082 -74798
rect 58150 -74804 58256 -74796
rect 58328 -74804 58434 -74796
rect 58508 -74804 58614 -74796
rect 58678 -74804 58784 -74796
rect 58858 -74804 58964 -74796
rect 59042 -74804 59148 -74796
rect 59216 -74804 59322 -74796
rect 59390 -74802 59496 -74796
rect 59568 -74798 59674 -74796
rect 59856 -74794 59926 -74642
rect 60032 -74794 60106 -74638
rect 60212 -74794 60278 -74638
rect 60384 -74642 60636 -74638
rect 60384 -74794 60462 -74642
rect 59856 -74796 60462 -74794
rect 59750 -74808 59856 -74798
rect 59926 -74804 60032 -74796
rect 60106 -74804 60212 -74796
rect 60278 -74804 60384 -74796
rect 60568 -74794 60636 -74642
rect 60742 -74642 61168 -74638
rect 60742 -74794 60816 -74642
rect 60568 -74796 60816 -74794
rect 60462 -74808 60568 -74798
rect 60636 -74804 60742 -74796
rect 60922 -74796 60992 -74642
rect 60816 -74808 60922 -74798
rect 61098 -74794 61168 -74642
rect 61274 -74642 61528 -74638
rect 61274 -74794 61348 -74642
rect 61098 -74796 61348 -74794
rect 60992 -74808 61098 -74798
rect 61168 -74804 61274 -74796
rect 61454 -74794 61528 -74642
rect 61634 -74646 61886 -74638
rect 61634 -74794 61706 -74646
rect 61454 -74796 61706 -74794
rect 61348 -74808 61454 -74798
rect 61528 -74804 61634 -74796
rect 61812 -74794 61886 -74646
rect 61992 -74642 62240 -74638
rect 61992 -74794 62062 -74642
rect 61812 -74796 62062 -74794
rect 61706 -74812 61812 -74802
rect 61886 -74804 61992 -74796
rect 62168 -74788 62240 -74642
rect 62346 -74636 64372 -74632
rect 62346 -74638 63848 -74636
rect 62346 -74788 62418 -74638
rect 62168 -74794 62418 -74788
rect 62524 -74794 62596 -74638
rect 62702 -74642 63130 -74638
rect 62702 -74794 62776 -74642
rect 62168 -74796 62776 -74794
rect 62240 -74798 62346 -74796
rect 62062 -74808 62168 -74798
rect 62418 -74804 62524 -74796
rect 62596 -74804 62702 -74796
rect 62882 -74796 62956 -74642
rect 62776 -74808 62882 -74798
rect 63062 -74794 63130 -74642
rect 63236 -74642 63848 -74638
rect 63236 -74794 63314 -74642
rect 63062 -74796 63314 -74794
rect 62956 -74808 63062 -74798
rect 63130 -74804 63236 -74796
rect 63420 -74796 63482 -74642
rect 63314 -74808 63420 -74798
rect 63588 -74648 63848 -74642
rect 63588 -74796 63660 -74648
rect 63482 -74808 63588 -74798
rect 63766 -74792 63848 -74648
rect 63954 -74638 64200 -74636
rect 63954 -74792 64020 -74638
rect 63766 -74794 64020 -74792
rect 64126 -74792 64200 -74638
rect 64306 -74792 64372 -74636
rect 64126 -74794 64306 -74792
rect 63766 -74796 64306 -74794
rect 63848 -74802 63954 -74796
rect 64020 -74804 64126 -74796
rect 64200 -74802 64306 -74796
rect 63660 -74814 63766 -74804
rect 56486 -74848 56520 -74840
rect 56842 -74848 56876 -74838
rect 56298 -74860 56352 -74850
rect 56474 -74854 56528 -74848
rect 56292 -76006 56298 -74861
rect 56292 -76016 56352 -76006
rect 56472 -74858 56528 -74854
rect 56652 -74855 56706 -74852
rect 56472 -74864 56474 -74858
rect 56472 -76004 56474 -76002
rect 56472 -76012 56528 -76004
rect 56474 -76014 56528 -76012
rect 56646 -74862 56706 -74855
rect 56646 -76008 56652 -74862
rect 56486 -76016 56520 -76014
rect 53804 -76772 54966 -76432
rect 56292 -76478 56346 -76016
rect 56646 -76018 56706 -76008
rect 56836 -74858 56892 -74848
rect 56890 -76004 56892 -75996
rect 56836 -76006 56892 -76004
rect 57010 -74866 57064 -74856
rect 57198 -74860 57232 -74838
rect 57554 -74852 57588 -74838
rect 57542 -74854 57596 -74852
rect 56836 -76014 56890 -76006
rect 57180 -74870 57240 -74860
rect 57064 -76012 57068 -74881
rect 56646 -76478 56700 -76018
rect 57010 -76022 57068 -76012
rect 57366 -74866 57420 -74856
rect 57180 -76016 57186 -76008
rect 57180 -76018 57240 -76016
rect 57014 -76478 57068 -76022
rect 57186 -76026 57240 -76018
rect 57360 -76012 57366 -74871
rect 57540 -74862 57596 -74854
rect 57540 -74864 57542 -74862
rect 57724 -74862 57778 -74852
rect 57908 -74856 57942 -74840
rect 57540 -76008 57542 -76002
rect 57540 -76012 57596 -76008
rect 57360 -76022 57420 -76012
rect 57542 -76018 57596 -76012
rect 57718 -76008 57724 -74871
rect 57718 -76018 57778 -76008
rect 57900 -74860 57954 -74856
rect 57900 -74866 57956 -74860
rect 57954 -74870 57956 -74866
rect 58078 -74866 58132 -74856
rect 58266 -74860 58300 -74838
rect 58622 -74852 58656 -74838
rect 58978 -74852 59012 -74840
rect 59334 -74852 59368 -74838
rect 58260 -74862 58314 -74860
rect 57954 -76012 57956 -76008
rect 57900 -76018 57956 -76012
rect 58072 -76012 58078 -74871
rect 57360 -76478 57414 -76022
rect 57718 -76478 57772 -76018
rect 57900 -76022 57954 -76018
rect 58072 -76022 58132 -76012
rect 58258 -74870 58314 -74862
rect 58258 -74872 58260 -74870
rect 58258 -76016 58260 -76010
rect 58258 -76020 58314 -76016
rect 58072 -76478 58126 -76022
rect 58260 -76026 58314 -76020
rect 58434 -74861 58488 -74856
rect 58434 -74866 58490 -74861
rect 58488 -76012 58490 -74866
rect 58612 -74862 58668 -74852
rect 58612 -76010 58614 -76000
rect 58434 -76022 58490 -76012
rect 58614 -76020 58668 -76010
rect 58790 -74855 58844 -74854
rect 58790 -74864 58848 -74855
rect 58970 -74856 59024 -74852
rect 58844 -76010 58848 -74864
rect 58790 -76020 58848 -76010
rect 58964 -74862 59024 -74856
rect 58964 -74866 58970 -74862
rect 58964 -76008 58970 -76004
rect 58964 -76014 59024 -76008
rect 58970 -76018 59024 -76014
rect 59150 -74862 59204 -74852
rect 58436 -76478 58490 -76022
rect 58794 -76478 58848 -76020
rect 59150 -76478 59204 -76008
rect 59326 -74862 59382 -74852
rect 59506 -74855 59560 -74848
rect 59690 -74852 59724 -74838
rect 59326 -76008 59328 -76000
rect 59326 -76010 59382 -76008
rect 59328 -76018 59382 -76010
rect 59496 -74858 59560 -74855
rect 59682 -74856 59736 -74852
rect 60046 -74856 60080 -74840
rect 59496 -76004 59506 -74858
rect 59496 -76014 59560 -76004
rect 59678 -74862 59736 -74856
rect 59860 -74861 59914 -74856
rect 59678 -74866 59682 -74862
rect 59678 -76008 59682 -76004
rect 59678 -76014 59736 -76008
rect 59496 -76478 59550 -76014
rect 59682 -76018 59736 -76014
rect 59858 -74866 59914 -74861
rect 60038 -74864 60092 -74856
rect 59858 -76012 59860 -74866
rect 59858 -76022 59914 -76012
rect 60036 -74866 60092 -74864
rect 60036 -74874 60038 -74866
rect 60036 -76022 60092 -76012
rect 60212 -74866 60266 -74856
rect 60402 -74860 60436 -74842
rect 60758 -74852 60792 -74842
rect 60752 -74858 60806 -74852
rect 61114 -74856 61148 -74842
rect 61470 -74854 61504 -74842
rect 61462 -74856 61516 -74854
rect 60390 -74862 60444 -74860
rect 60572 -74861 60626 -74860
rect 60386 -74870 60444 -74862
rect 60266 -76012 60270 -74871
rect 60212 -76022 60270 -76012
rect 60386 -74872 60390 -74870
rect 60386 -76016 60390 -76010
rect 60386 -76020 60444 -76016
rect 59858 -76478 59912 -76022
rect 60216 -76478 60270 -76022
rect 60390 -76026 60444 -76020
rect 60562 -74870 60626 -74861
rect 60562 -76016 60572 -74870
rect 60748 -74862 60806 -74858
rect 60928 -74861 60982 -74856
rect 60748 -74868 60752 -74862
rect 60748 -76008 60752 -76006
rect 60748 -76016 60806 -76008
rect 60562 -76026 60626 -76016
rect 60752 -76018 60806 -76016
rect 60926 -74866 60982 -74861
rect 61106 -74862 61160 -74856
rect 61282 -74861 61336 -74860
rect 60926 -76012 60928 -74866
rect 60926 -76022 60982 -76012
rect 61102 -74866 61160 -74862
rect 61102 -74872 61106 -74866
rect 61102 -76012 61106 -76010
rect 61102 -76020 61160 -76012
rect 61106 -76022 61160 -76020
rect 61276 -74870 61336 -74861
rect 61276 -76016 61282 -74870
rect 61460 -74864 61516 -74856
rect 61460 -74866 61462 -74864
rect 61640 -74862 61694 -74852
rect 61826 -74856 61860 -74844
rect 62182 -74856 62216 -74846
rect 62538 -74854 62572 -74842
rect 61812 -74862 61866 -74856
rect 61460 -76010 61462 -76004
rect 61460 -76014 61516 -76010
rect 60562 -76478 60616 -76026
rect 60926 -76478 60980 -76022
rect 61276 -76026 61336 -76016
rect 61462 -76020 61516 -76014
rect 61634 -76008 61640 -74881
rect 61634 -76018 61694 -76008
rect 61810 -74866 61866 -74862
rect 61810 -74872 61812 -74866
rect 61810 -76012 61812 -76010
rect 61276 -76478 61330 -76026
rect 61634 -76478 61688 -76018
rect 61810 -76020 61866 -76012
rect 61812 -76022 61866 -76020
rect 61992 -74866 62046 -74856
rect 62172 -74866 62226 -74856
rect 62352 -74861 62406 -74856
rect 62340 -74866 62406 -74861
rect 62530 -74862 62584 -74854
rect 62226 -74876 62228 -74866
rect 62046 -76012 62048 -74881
rect 61992 -76022 62048 -76012
rect 61994 -76478 62048 -76022
rect 62172 -76024 62228 -76014
rect 62340 -76012 62352 -74866
rect 62340 -76022 62406 -76012
rect 62528 -74864 62584 -74862
rect 62528 -74872 62530 -74864
rect 62528 -76020 62584 -76010
rect 62704 -74860 62758 -74850
rect 62894 -74856 62928 -74840
rect 63250 -74850 63284 -74840
rect 62758 -76006 62760 -74861
rect 62882 -74866 62936 -74856
rect 62704 -76016 62760 -76006
rect 62340 -76478 62394 -76022
rect 62706 -76478 62760 -76016
rect 62878 -74876 62882 -74866
rect 63064 -74864 63118 -74854
rect 63240 -74860 63294 -74850
rect 63606 -74852 63640 -74840
rect 63962 -74850 63996 -74840
rect 62934 -76014 62936 -76012
rect 62878 -76022 62936 -76014
rect 63062 -76010 63064 -74881
rect 63062 -76020 63118 -76010
rect 63238 -74874 63240 -74864
rect 63416 -74864 63470 -74854
rect 62878 -76024 62934 -76022
rect 63062 -76478 63116 -76020
rect 63238 -76022 63294 -76012
rect 63412 -76010 63416 -74871
rect 63412 -76020 63470 -76010
rect 63596 -74862 63650 -74852
rect 63774 -74862 63828 -74852
rect 63952 -74860 64006 -74850
rect 63650 -74876 63654 -74866
rect 63596 -76014 63598 -76008
rect 63596 -76018 63654 -76014
rect 63412 -76478 63466 -76020
rect 63598 -76024 63654 -76018
rect 63770 -76008 63774 -74871
rect 63770 -76018 63828 -76008
rect 63950 -74870 63952 -74860
rect 63950 -76018 64006 -76008
rect 64130 -74858 64184 -74848
rect 64318 -74852 64352 -74842
rect 64306 -74860 64360 -74852
rect 63770 -76478 63824 -76018
rect 64130 -76478 64184 -76004
rect 64304 -74862 64360 -74860
rect 64304 -74870 64306 -74862
rect 64304 -76018 64360 -76008
rect 64468 -76478 66630 -73154
rect 67974 -73358 86894 -72930
rect 67974 -73360 84819 -73358
rect 56226 -76752 66630 -76478
rect 54815 -78492 54962 -76772
rect 56300 -77238 56354 -76752
rect 56492 -77236 56526 -77228
rect 56300 -77248 56358 -77238
rect 56480 -77242 56534 -77236
rect 56300 -78394 56304 -77248
rect 56300 -78403 56358 -78394
rect 56478 -77246 56534 -77242
rect 56478 -77252 56480 -77246
rect 56478 -78392 56480 -78390
rect 56478 -78400 56534 -78392
rect 56654 -77240 56708 -76752
rect 56848 -77236 56882 -77226
rect 56654 -77250 56712 -77240
rect 56654 -78393 56658 -77250
rect 56480 -78402 56534 -78400
rect 56304 -78404 56358 -78403
rect 56492 -78404 56526 -78402
rect 56658 -78406 56712 -78396
rect 56842 -77246 56898 -77236
rect 56896 -78392 56898 -78384
rect 56842 -78394 56898 -78392
rect 57010 -77244 57064 -76752
rect 57010 -77254 57070 -77244
rect 57204 -77248 57238 -77226
rect 57368 -77244 57422 -76752
rect 57560 -77240 57594 -77226
rect 57718 -77240 57772 -76752
rect 57548 -77242 57602 -77240
rect 56842 -78402 56896 -78394
rect 57010 -78400 57016 -77254
rect 57010 -78409 57070 -78400
rect 57186 -77258 57246 -77248
rect 57186 -78404 57192 -78396
rect 57186 -78406 57246 -78404
rect 57016 -78410 57070 -78409
rect 57192 -78414 57246 -78406
rect 57368 -77254 57426 -77244
rect 57368 -78400 57372 -77254
rect 57546 -77250 57602 -77242
rect 57546 -77252 57548 -77250
rect 57546 -78396 57548 -78390
rect 57546 -78400 57602 -78396
rect 57368 -78410 57426 -78400
rect 57548 -78406 57602 -78400
rect 57718 -77250 57784 -77240
rect 57914 -77244 57948 -77228
rect 58082 -77244 58136 -76752
rect 57718 -78396 57730 -77250
rect 57718 -78406 57784 -78396
rect 57906 -77248 57960 -77244
rect 57906 -77254 57962 -77248
rect 57960 -77258 57962 -77254
rect 57960 -78400 57962 -78396
rect 57906 -78406 57962 -78400
rect 58082 -77254 58138 -77244
rect 58272 -77248 58306 -77226
rect 58432 -77244 58486 -76752
rect 58628 -77240 58662 -77226
rect 58266 -77250 58320 -77248
rect 58082 -78400 58084 -77254
rect 58082 -78403 58138 -78400
rect 57718 -78409 57772 -78406
rect 57906 -78410 57960 -78406
rect 58084 -78410 58138 -78403
rect 58264 -77258 58320 -77250
rect 58264 -77260 58266 -77258
rect 58264 -78404 58266 -78398
rect 58264 -78408 58320 -78404
rect 57368 -78419 57422 -78410
rect 58266 -78414 58320 -78408
rect 58432 -77254 58494 -77244
rect 58432 -78400 58440 -77254
rect 58618 -77250 58674 -77240
rect 58618 -78398 58620 -78388
rect 58790 -77242 58844 -76752
rect 58984 -77240 59018 -77228
rect 59146 -77240 59200 -76752
rect 59340 -77240 59374 -77226
rect 59496 -77236 59550 -76752
rect 58790 -77252 58850 -77242
rect 58976 -77244 59030 -77240
rect 58790 -78393 58796 -77252
rect 58432 -78409 58494 -78400
rect 58620 -78408 58674 -78398
rect 58796 -78408 58850 -78398
rect 58970 -77250 59030 -77244
rect 58970 -77254 58976 -77250
rect 58970 -78396 58976 -78392
rect 59146 -77250 59210 -77240
rect 59146 -78393 59156 -77250
rect 58970 -78402 59030 -78396
rect 58976 -78406 59030 -78402
rect 59156 -78406 59210 -78396
rect 59332 -77250 59388 -77240
rect 59332 -78396 59334 -78388
rect 59332 -78398 59388 -78396
rect 59334 -78406 59388 -78398
rect 59496 -77246 59566 -77236
rect 59696 -77240 59730 -77226
rect 59688 -77244 59742 -77240
rect 59870 -77244 59924 -76752
rect 60052 -77244 60086 -77228
rect 60216 -77244 60270 -76752
rect 59496 -78392 59512 -77246
rect 59496 -78402 59566 -78392
rect 59684 -77250 59742 -77244
rect 59684 -77254 59688 -77250
rect 59684 -78396 59688 -78392
rect 59684 -78402 59742 -78396
rect 59496 -78403 59550 -78402
rect 59688 -78406 59742 -78402
rect 59866 -77254 59924 -77244
rect 60044 -77252 60098 -77244
rect 59920 -78400 59924 -77254
rect 58440 -78410 58494 -78409
rect 59866 -78409 59924 -78400
rect 60042 -77254 60098 -77252
rect 60042 -77262 60044 -77254
rect 59866 -78410 59920 -78409
rect 60042 -78410 60098 -78400
rect 60216 -77254 60272 -77244
rect 60408 -77248 60442 -77230
rect 60576 -77248 60630 -76752
rect 60764 -77240 60798 -77230
rect 60758 -77246 60812 -77240
rect 60396 -77250 60450 -77248
rect 60216 -78400 60218 -77254
rect 60216 -78409 60272 -78400
rect 60392 -77258 60450 -77250
rect 60392 -77260 60396 -77258
rect 60392 -78404 60396 -78398
rect 60392 -78408 60450 -78404
rect 60218 -78410 60272 -78409
rect 60396 -78414 60450 -78408
rect 60576 -77258 60632 -77248
rect 60576 -78404 60578 -77258
rect 60754 -77250 60812 -77246
rect 60754 -77256 60758 -77250
rect 60754 -78396 60758 -78394
rect 60754 -78404 60812 -78396
rect 60576 -78409 60632 -78404
rect 60758 -78406 60812 -78404
rect 60934 -77254 60988 -76752
rect 61120 -77244 61154 -77230
rect 61112 -77250 61166 -77244
rect 60578 -78414 60632 -78409
rect 60934 -78410 60988 -78400
rect 61108 -77254 61166 -77250
rect 61108 -77260 61112 -77254
rect 61108 -78400 61112 -78398
rect 61108 -78408 61166 -78400
rect 61112 -78410 61166 -78408
rect 61288 -77258 61342 -76752
rect 61476 -77242 61510 -77230
rect 61644 -77240 61698 -76752
rect 61468 -77244 61522 -77242
rect 61466 -77252 61522 -77244
rect 61466 -77254 61468 -77252
rect 61466 -78398 61468 -78392
rect 61466 -78402 61522 -78398
rect 61288 -78414 61342 -78404
rect 61468 -78408 61522 -78402
rect 61644 -77250 61700 -77240
rect 61832 -77244 61866 -77232
rect 62002 -77244 62056 -76752
rect 62188 -77244 62222 -77234
rect 62360 -77244 62414 -76752
rect 62544 -77242 62578 -77230
rect 62716 -77238 62770 -76752
rect 61818 -77250 61872 -77244
rect 61644 -78396 61646 -77250
rect 61644 -78403 61700 -78396
rect 61646 -78406 61700 -78403
rect 61816 -77254 61872 -77250
rect 61816 -77260 61818 -77254
rect 61816 -78400 61818 -78398
rect 61816 -78408 61872 -78400
rect 61818 -78410 61872 -78408
rect 61998 -77254 62056 -77244
rect 62052 -78400 62056 -77254
rect 61998 -78410 62056 -78400
rect 62002 -78419 62056 -78410
rect 62178 -77254 62232 -77244
rect 62358 -77254 62414 -77244
rect 62536 -77250 62590 -77242
rect 62232 -77264 62234 -77254
rect 62178 -78412 62234 -78402
rect 62412 -78400 62414 -77254
rect 62358 -78410 62414 -78400
rect 62534 -77252 62590 -77250
rect 62534 -77260 62536 -77252
rect 62534 -78408 62590 -78398
rect 62710 -77248 62770 -77238
rect 62900 -77244 62934 -77228
rect 63066 -77242 63120 -76752
rect 63256 -77238 63290 -77228
rect 62764 -78394 62770 -77248
rect 62888 -77254 62942 -77244
rect 62710 -78404 62770 -78394
rect 62360 -78419 62414 -78410
rect 62716 -78425 62770 -78404
rect 62884 -77264 62888 -77254
rect 62940 -78402 62942 -78400
rect 62884 -78410 62942 -78402
rect 63066 -77252 63124 -77242
rect 63246 -77248 63300 -77238
rect 63424 -77242 63478 -76752
rect 63612 -77240 63646 -77228
rect 63782 -77240 63836 -76752
rect 63968 -77238 64002 -77228
rect 64134 -77236 64188 -76752
rect 63066 -78398 63070 -77252
rect 63066 -78408 63124 -78398
rect 63244 -77262 63246 -77252
rect 63066 -78409 63120 -78408
rect 63244 -78410 63300 -78400
rect 63422 -77252 63478 -77242
rect 63476 -78393 63478 -77252
rect 63602 -77250 63656 -77240
rect 63780 -77250 63836 -77240
rect 63958 -77248 64012 -77238
rect 63656 -77264 63660 -77254
rect 63422 -78408 63476 -78398
rect 63602 -78402 63604 -78396
rect 63602 -78406 63660 -78402
rect 63834 -78396 63836 -77250
rect 63780 -78406 63836 -78396
rect 63956 -77258 63958 -77248
rect 64134 -77246 64190 -77236
rect 64324 -77240 64358 -77230
rect 64134 -78392 64136 -77246
rect 64312 -77248 64366 -77240
rect 64134 -78393 64190 -78392
rect 63956 -78406 64012 -78396
rect 64136 -78402 64190 -78393
rect 64310 -77250 64366 -77248
rect 64310 -77258 64312 -77250
rect 64310 -78406 64366 -78396
rect 62884 -78412 62940 -78410
rect 63604 -78412 63660 -78406
rect 63782 -78419 63836 -78406
rect 56354 -78486 56460 -78476
rect 54814 -78642 56354 -78492
rect 56536 -78492 56642 -78482
rect 56718 -78488 56824 -78478
rect 56460 -78642 56536 -78492
rect 54814 -78648 56536 -78642
rect 56642 -78644 56718 -78492
rect 56898 -78488 57004 -78478
rect 56824 -78644 56898 -78492
rect 57076 -78486 57182 -78476
rect 57004 -78642 57076 -78492
rect 57252 -78486 57358 -78476
rect 57182 -78642 57252 -78492
rect 57436 -78488 57542 -78478
rect 57358 -78642 57436 -78492
rect 57004 -78644 57436 -78642
rect 57610 -78488 57716 -78478
rect 57542 -78644 57610 -78492
rect 57784 -78488 57890 -78478
rect 57716 -78644 57784 -78492
rect 57966 -78492 58072 -78482
rect 58140 -78488 58246 -78478
rect 57890 -78644 57966 -78492
rect 56642 -78648 57966 -78644
rect 58072 -78644 58140 -78492
rect 58318 -78488 58424 -78478
rect 58246 -78644 58318 -78492
rect 58498 -78488 58604 -78478
rect 58424 -78644 58498 -78492
rect 58668 -78488 58774 -78478
rect 58604 -78644 58668 -78492
rect 58848 -78488 58954 -78478
rect 58774 -78644 58848 -78492
rect 59032 -78488 59138 -78478
rect 58954 -78644 59032 -78492
rect 59206 -78488 59312 -78478
rect 59138 -78644 59206 -78492
rect 59380 -78486 59486 -78476
rect 59312 -78642 59380 -78492
rect 59558 -78482 59664 -78472
rect 59486 -78638 59558 -78492
rect 59740 -78492 59846 -78482
rect 59916 -78488 60022 -78478
rect 59664 -78638 59740 -78492
rect 59486 -78642 59740 -78638
rect 59312 -78644 59740 -78642
rect 58072 -78648 59740 -78644
rect 59846 -78644 59916 -78492
rect 60096 -78488 60202 -78478
rect 60022 -78644 60096 -78492
rect 60268 -78488 60374 -78478
rect 60202 -78644 60268 -78492
rect 60452 -78492 60558 -78482
rect 60626 -78488 60732 -78478
rect 60374 -78644 60452 -78492
rect 59846 -78648 60452 -78644
rect 60558 -78644 60626 -78492
rect 60806 -78492 60912 -78482
rect 60982 -78492 61088 -78482
rect 61158 -78488 61264 -78478
rect 60732 -78644 60806 -78492
rect 60558 -78648 60806 -78644
rect 60912 -78648 60982 -78492
rect 61088 -78644 61158 -78492
rect 61338 -78492 61444 -78482
rect 61518 -78488 61624 -78478
rect 61264 -78644 61338 -78492
rect 61088 -78648 61338 -78644
rect 61444 -78644 61518 -78492
rect 61696 -78492 61802 -78486
rect 61876 -78488 61982 -78478
rect 62230 -78482 62336 -78472
rect 61624 -78496 61876 -78492
rect 61624 -78644 61696 -78496
rect 61444 -78648 61696 -78644
rect 54814 -78652 61696 -78648
rect 61802 -78644 61876 -78496
rect 62052 -78492 62158 -78482
rect 61982 -78644 62052 -78492
rect 61802 -78648 62052 -78644
rect 62158 -78638 62230 -78492
rect 62408 -78488 62514 -78478
rect 62336 -78638 62408 -78492
rect 62158 -78644 62408 -78638
rect 62586 -78488 62692 -78478
rect 62514 -78644 62586 -78492
rect 62766 -78492 62872 -78482
rect 62946 -78492 63052 -78482
rect 63120 -78488 63226 -78478
rect 62692 -78644 62766 -78492
rect 62158 -78648 62766 -78644
rect 62872 -78648 62946 -78492
rect 63052 -78644 63120 -78492
rect 63304 -78492 63410 -78482
rect 63472 -78492 63578 -78482
rect 63838 -78486 63944 -78476
rect 63650 -78492 63756 -78488
rect 63226 -78644 63304 -78492
rect 63052 -78648 63304 -78644
rect 63410 -78648 63472 -78492
rect 63578 -78498 63838 -78492
rect 63578 -78648 63650 -78498
rect 61802 -78652 63650 -78648
rect 54814 -78654 63650 -78652
rect 63756 -78642 63838 -78498
rect 64010 -78488 64116 -78478
rect 63944 -78642 64010 -78492
rect 63756 -78644 64010 -78642
rect 64190 -78486 64296 -78476
rect 64116 -78642 64190 -78492
rect 64296 -78494 64306 -78492
rect 64296 -78642 64366 -78494
rect 64116 -78644 64366 -78642
rect 63756 -78654 64366 -78644
rect 54814 -78658 64366 -78654
rect 61696 -78662 61802 -78658
rect 63650 -78664 63756 -78658
rect 56292 -78700 56346 -78689
rect 56476 -78698 56510 -78690
rect 56832 -78698 56866 -78688
rect 56288 -78710 56346 -78700
rect 56464 -78704 56518 -78698
rect 56342 -79856 56346 -78710
rect 56288 -79866 56346 -79856
rect 56462 -78708 56518 -78704
rect 56462 -78714 56464 -78708
rect 56462 -79854 56464 -79852
rect 56462 -79862 56518 -79854
rect 56464 -79864 56518 -79862
rect 56642 -78712 56696 -78702
rect 56826 -78708 56882 -78698
rect 56696 -79858 56700 -78715
rect 56476 -79866 56510 -79864
rect 56292 -80470 56346 -79866
rect 56642 -79868 56700 -79858
rect 56880 -79854 56882 -79846
rect 56826 -79856 56882 -79854
rect 57000 -78716 57054 -78706
rect 57188 -78710 57222 -78688
rect 57544 -78702 57578 -78688
rect 57532 -78704 57586 -78702
rect 56826 -79864 56880 -79856
rect 57170 -78720 57230 -78710
rect 57054 -79862 57068 -78725
rect 56646 -80470 56700 -79868
rect 57000 -79872 57068 -79862
rect 57170 -79866 57176 -79858
rect 57170 -79868 57230 -79866
rect 57014 -80470 57068 -79872
rect 57176 -79876 57230 -79868
rect 57356 -78716 57410 -78706
rect 57530 -78712 57586 -78704
rect 57530 -78714 57532 -78712
rect 57410 -79862 57414 -78725
rect 57530 -79858 57532 -79852
rect 57530 -79862 57586 -79858
rect 57356 -79872 57414 -79862
rect 57532 -79868 57586 -79862
rect 57714 -78712 57768 -78702
rect 57898 -78706 57932 -78690
rect 57890 -78710 57944 -78706
rect 57890 -78716 57946 -78710
rect 57944 -78720 57946 -78716
rect 57768 -79858 57772 -78725
rect 57714 -79868 57772 -79858
rect 57360 -80470 57414 -79872
rect 57718 -80470 57772 -79868
rect 57944 -79862 57946 -79858
rect 57890 -79868 57946 -79862
rect 58068 -78716 58122 -78706
rect 58256 -78710 58290 -78688
rect 58612 -78702 58646 -78688
rect 58968 -78702 59002 -78690
rect 59324 -78702 59358 -78688
rect 58250 -78712 58304 -78710
rect 58248 -78720 58304 -78712
rect 58248 -78722 58250 -78720
rect 58122 -79862 58126 -78731
rect 57890 -79872 57944 -79868
rect 58068 -79872 58126 -79862
rect 58248 -79866 58250 -79860
rect 58248 -79870 58304 -79866
rect 58072 -80470 58126 -79872
rect 58250 -79876 58304 -79870
rect 58424 -78716 58478 -78706
rect 58602 -78712 58658 -78702
rect 58478 -79862 58490 -78731
rect 58602 -79860 58604 -79850
rect 58424 -79872 58490 -79862
rect 58604 -79870 58658 -79860
rect 58780 -78714 58834 -78704
rect 58960 -78706 59014 -78702
rect 58954 -78712 59014 -78706
rect 58954 -78716 58960 -78712
rect 58834 -79860 58848 -78725
rect 58780 -79870 58848 -79860
rect 58954 -79858 58960 -79854
rect 58954 -79864 59014 -79858
rect 58960 -79868 59014 -79864
rect 59140 -78709 59194 -78702
rect 59140 -78712 59204 -78709
rect 59194 -79858 59204 -78712
rect 59140 -79868 59204 -79858
rect 59316 -78712 59372 -78702
rect 59316 -79858 59318 -79850
rect 59316 -79860 59372 -79858
rect 59318 -79868 59372 -79860
rect 59496 -78708 59550 -78698
rect 59680 -78702 59714 -78688
rect 59672 -78706 59726 -78702
rect 59866 -78706 59920 -78689
rect 60036 -78706 60070 -78690
rect 58436 -80470 58490 -79872
rect 58794 -80470 58848 -79870
rect 59150 -80470 59204 -79868
rect 59496 -80470 59550 -79854
rect 59668 -78712 59726 -78706
rect 59668 -78716 59672 -78712
rect 59668 -79858 59672 -79854
rect 59668 -79864 59726 -79858
rect 59672 -79868 59726 -79864
rect 59850 -78716 59920 -78706
rect 60028 -78714 60082 -78706
rect 59904 -79862 59920 -78716
rect 59850 -79872 59920 -79862
rect 60026 -78716 60082 -78714
rect 60026 -78724 60028 -78716
rect 60026 -79872 60082 -79862
rect 60202 -78716 60256 -78706
rect 60392 -78710 60426 -78692
rect 60748 -78702 60782 -78692
rect 60742 -78708 60796 -78702
rect 61104 -78706 61138 -78692
rect 60380 -78712 60434 -78710
rect 60376 -78720 60434 -78712
rect 60376 -78722 60380 -78720
rect 60256 -79862 60278 -78725
rect 60202 -79872 60278 -79862
rect 60376 -79866 60380 -79860
rect 60376 -79870 60434 -79866
rect 59866 -80470 59920 -79872
rect 60224 -80470 60278 -79872
rect 60380 -79876 60434 -79870
rect 60562 -78720 60616 -78710
rect 60738 -78712 60796 -78708
rect 60738 -78718 60742 -78712
rect 60616 -79866 60624 -78725
rect 60738 -79858 60742 -79856
rect 60738 -79866 60796 -79858
rect 60562 -79876 60624 -79866
rect 60742 -79868 60796 -79866
rect 60918 -78715 60972 -78706
rect 61096 -78712 61150 -78706
rect 61284 -78710 61338 -78699
rect 61460 -78704 61494 -78692
rect 61452 -78706 61506 -78704
rect 60918 -78716 60988 -78715
rect 60972 -79862 60988 -78716
rect 60918 -79872 60988 -79862
rect 61092 -78716 61150 -78712
rect 61092 -78722 61096 -78716
rect 61092 -79862 61096 -79860
rect 61092 -79870 61150 -79862
rect 61096 -79872 61150 -79870
rect 61272 -78720 61338 -78710
rect 61326 -79866 61338 -78720
rect 61450 -78714 61506 -78706
rect 61450 -78716 61452 -78714
rect 61450 -79860 61452 -79854
rect 61450 -79864 61506 -79860
rect 60570 -80470 60624 -79876
rect 60934 -80470 60988 -79872
rect 61272 -79876 61338 -79866
rect 61452 -79870 61506 -79864
rect 61630 -78712 61684 -78702
rect 61816 -78706 61850 -78694
rect 62172 -78706 62206 -78696
rect 62528 -78704 62562 -78692
rect 61802 -78712 61856 -78706
rect 61800 -78716 61856 -78712
rect 61800 -78722 61802 -78716
rect 61684 -79858 61696 -78725
rect 61630 -79868 61696 -79858
rect 61284 -80470 61338 -79876
rect 61642 -80470 61696 -79868
rect 61800 -79862 61802 -79860
rect 61800 -79870 61856 -79862
rect 61802 -79872 61856 -79870
rect 61982 -78709 62036 -78706
rect 61982 -78716 62056 -78709
rect 62036 -79862 62056 -78716
rect 61982 -79872 62056 -79862
rect 62002 -80470 62056 -79872
rect 62162 -78716 62216 -78706
rect 62342 -78716 62396 -78706
rect 62520 -78712 62574 -78704
rect 62216 -78726 62218 -78716
rect 62162 -79874 62218 -79864
rect 62518 -78714 62574 -78712
rect 62518 -78722 62520 -78714
rect 62396 -79862 62402 -78731
rect 62342 -79872 62402 -79862
rect 62518 -79870 62574 -79860
rect 62694 -78710 62748 -78700
rect 62884 -78706 62918 -78690
rect 63240 -78700 63274 -78690
rect 62748 -79856 62768 -78715
rect 62872 -78716 62926 -78706
rect 62694 -79866 62768 -79856
rect 62348 -80470 62402 -79872
rect 62714 -80470 62768 -79866
rect 62868 -78726 62872 -78716
rect 62924 -79864 62926 -79862
rect 62868 -79872 62926 -79864
rect 63054 -78714 63108 -78704
rect 63230 -78710 63284 -78700
rect 63596 -78702 63630 -78690
rect 63952 -78700 63986 -78690
rect 63108 -79860 63124 -78715
rect 63054 -79870 63124 -79860
rect 62868 -79874 62924 -79872
rect 63070 -80470 63124 -79870
rect 63228 -78724 63230 -78714
rect 63228 -79872 63284 -79862
rect 63406 -78714 63460 -78704
rect 63586 -78712 63640 -78702
rect 63460 -79860 63474 -78715
rect 63406 -79870 63474 -79860
rect 63764 -78712 63818 -78702
rect 63942 -78710 63996 -78700
rect 63640 -78726 63644 -78716
rect 63586 -79864 63588 -79858
rect 63586 -79868 63644 -79864
rect 63818 -79858 63832 -78715
rect 63764 -79868 63832 -79858
rect 63940 -78720 63942 -78710
rect 63940 -79868 63996 -79858
rect 64120 -78708 64174 -78698
rect 64308 -78702 64342 -78692
rect 64174 -79854 64192 -78709
rect 64296 -78710 64350 -78702
rect 64120 -79864 64192 -79854
rect 63420 -80470 63474 -79870
rect 63588 -79874 63644 -79868
rect 63778 -80470 63832 -79868
rect 64138 -80470 64192 -79864
rect 64294 -78712 64350 -78710
rect 64294 -78720 64296 -78712
rect 64294 -79868 64350 -79858
rect 64468 -80470 66630 -76752
rect 56199 -80744 66630 -80470
rect 56298 -81204 56352 -80744
rect 56502 -81202 56536 -81194
rect 56298 -81214 56368 -81204
rect 56490 -81208 56544 -81202
rect 56298 -82360 56314 -81214
rect 56298 -82365 56368 -82360
rect 56314 -82370 56368 -82365
rect 56488 -81212 56544 -81208
rect 56488 -81218 56490 -81212
rect 56488 -82358 56490 -82356
rect 56488 -82366 56544 -82358
rect 56490 -82368 56544 -82366
rect 56652 -81206 56706 -80744
rect 56858 -81202 56892 -81192
rect 56652 -81216 56722 -81206
rect 56652 -82362 56668 -81216
rect 56502 -82370 56536 -82368
rect 56652 -82372 56722 -82362
rect 56852 -81212 56908 -81202
rect 56906 -82358 56908 -82350
rect 56852 -82360 56908 -82358
rect 57008 -81210 57062 -80744
rect 57008 -81220 57080 -81210
rect 57214 -81214 57248 -81192
rect 57366 -81210 57420 -80744
rect 57570 -81206 57604 -81192
rect 57716 -81206 57770 -80744
rect 57558 -81208 57612 -81206
rect 56852 -82368 56906 -82360
rect 57008 -82366 57026 -81220
rect 57008 -82371 57080 -82366
rect 56652 -82403 56706 -82372
rect 57026 -82376 57080 -82371
rect 57196 -81224 57256 -81214
rect 57366 -81220 57436 -81210
rect 57366 -82355 57382 -81220
rect 57196 -82370 57202 -82362
rect 57196 -82372 57256 -82370
rect 57202 -82380 57256 -82372
rect 57556 -81216 57612 -81208
rect 57556 -81218 57558 -81216
rect 57556 -82362 57558 -82356
rect 57556 -82366 57612 -82362
rect 57382 -82376 57436 -82366
rect 57558 -82372 57612 -82366
rect 57716 -81216 57794 -81206
rect 57924 -81210 57958 -81194
rect 58080 -81210 58134 -80744
rect 57716 -82362 57740 -81216
rect 57716 -82371 57794 -82362
rect 57740 -82372 57794 -82371
rect 57916 -81214 57970 -81210
rect 57916 -81220 57972 -81214
rect 57970 -81224 57972 -81220
rect 58080 -81220 58148 -81210
rect 58282 -81214 58316 -81192
rect 58430 -81210 58484 -80744
rect 58638 -81206 58672 -81192
rect 58276 -81216 58330 -81214
rect 58080 -82361 58094 -81220
rect 57970 -82366 57972 -82362
rect 57916 -82372 57972 -82366
rect 57916 -82376 57970 -82372
rect 58094 -82376 58148 -82366
rect 58274 -81224 58330 -81216
rect 58274 -81226 58276 -81224
rect 58274 -82370 58276 -82364
rect 58274 -82374 58330 -82370
rect 58276 -82380 58330 -82374
rect 58430 -81220 58504 -81210
rect 58430 -82366 58450 -81220
rect 58628 -81216 58684 -81206
rect 58628 -82364 58630 -82354
rect 58430 -82376 58504 -82366
rect 58630 -82374 58684 -82364
rect 58788 -81208 58842 -80744
rect 58994 -81206 59028 -81194
rect 59144 -81206 59198 -80744
rect 59350 -81206 59384 -81192
rect 59494 -81202 59548 -80744
rect 58788 -81218 58860 -81208
rect 58986 -81210 59040 -81206
rect 58788 -82364 58806 -81218
rect 58788 -82371 58860 -82364
rect 58980 -81216 59040 -81210
rect 58980 -81220 58986 -81216
rect 58980 -82362 58986 -82358
rect 58980 -82368 59040 -82362
rect 58806 -82374 58860 -82371
rect 58986 -82372 59040 -82368
rect 59144 -81216 59220 -81206
rect 59144 -82362 59166 -81216
rect 59144 -82371 59220 -82362
rect 59342 -81216 59398 -81206
rect 59342 -82362 59344 -82354
rect 59342 -82364 59398 -82362
rect 59166 -82372 59220 -82371
rect 59344 -82372 59398 -82364
rect 59494 -81212 59576 -81202
rect 59706 -81206 59740 -81192
rect 59698 -81210 59752 -81206
rect 59494 -82358 59522 -81212
rect 59494 -82368 59576 -82358
rect 59694 -81216 59752 -81210
rect 59694 -81220 59698 -81216
rect 59694 -82362 59698 -82358
rect 59694 -82368 59752 -82362
rect 58430 -82387 58484 -82376
rect 59494 -82383 59548 -82368
rect 59698 -82372 59752 -82368
rect 59860 -81210 59914 -80744
rect 60062 -81210 60096 -81194
rect 60206 -81210 60260 -80744
rect 59860 -81220 59930 -81210
rect 60054 -81218 60108 -81210
rect 59860 -82366 59876 -81220
rect 59860 -82376 59930 -82366
rect 60052 -81220 60108 -81218
rect 60052 -81228 60054 -81220
rect 60052 -82376 60108 -82366
rect 60206 -81220 60282 -81210
rect 60418 -81214 60452 -81196
rect 60566 -81214 60620 -80744
rect 60774 -81206 60808 -81196
rect 60768 -81212 60822 -81206
rect 60406 -81216 60460 -81214
rect 60206 -82366 60228 -81220
rect 60206 -82371 60282 -82366
rect 60228 -82376 60282 -82371
rect 60402 -81224 60460 -81216
rect 60402 -81226 60406 -81224
rect 60402 -82370 60406 -82364
rect 60402 -82374 60460 -82370
rect 59860 -82387 59914 -82376
rect 60406 -82380 60460 -82374
rect 60566 -81224 60642 -81214
rect 60566 -82370 60588 -81224
rect 60764 -81216 60822 -81212
rect 60764 -81222 60768 -81216
rect 60764 -82362 60768 -82360
rect 60764 -82370 60822 -82362
rect 60566 -82380 60642 -82370
rect 60768 -82372 60822 -82370
rect 60924 -81210 60978 -80744
rect 61130 -81210 61164 -81196
rect 60924 -81220 60998 -81210
rect 61122 -81216 61176 -81210
rect 60924 -82366 60944 -81220
rect 60924 -82376 60998 -82366
rect 61118 -81220 61176 -81216
rect 61118 -81226 61122 -81220
rect 61118 -82366 61122 -82364
rect 61118 -82374 61176 -82366
rect 61278 -81214 61332 -80744
rect 61486 -81208 61520 -81196
rect 61634 -81206 61688 -80744
rect 61478 -81210 61532 -81208
rect 61278 -81224 61352 -81214
rect 61278 -82370 61298 -81224
rect 61476 -81218 61532 -81210
rect 61476 -81220 61478 -81218
rect 61476 -82364 61478 -82358
rect 61476 -82368 61532 -82364
rect 61278 -82371 61352 -82370
rect 61122 -82376 61176 -82374
rect 60566 -82387 60620 -82380
rect 60924 -82399 60978 -82376
rect 61298 -82380 61352 -82371
rect 61478 -82374 61532 -82368
rect 61634 -81216 61710 -81206
rect 61842 -81210 61876 -81198
rect 61992 -81210 62046 -80744
rect 62198 -81210 62232 -81200
rect 62350 -81210 62404 -80744
rect 62554 -81208 62588 -81196
rect 62706 -81204 62760 -80744
rect 61828 -81216 61882 -81210
rect 61634 -82362 61656 -81216
rect 61634 -82371 61710 -82362
rect 61656 -82372 61710 -82371
rect 61826 -81220 61882 -81216
rect 61826 -81226 61828 -81220
rect 61826 -82366 61828 -82364
rect 61826 -82374 61882 -82366
rect 61992 -81220 62062 -81210
rect 61992 -82366 62008 -81220
rect 61992 -82371 62062 -82366
rect 61828 -82376 61882 -82374
rect 62008 -82376 62062 -82371
rect 62188 -81220 62242 -81210
rect 62350 -81220 62422 -81210
rect 62546 -81216 62600 -81208
rect 62242 -81230 62244 -81220
rect 62188 -82378 62244 -82368
rect 62350 -82366 62368 -81220
rect 62350 -82376 62422 -82366
rect 62544 -81218 62600 -81216
rect 62544 -81226 62546 -81218
rect 62706 -81214 62774 -81204
rect 62910 -81210 62944 -81194
rect 63056 -81208 63110 -80744
rect 63266 -81204 63300 -81194
rect 62706 -82360 62720 -81214
rect 62898 -81220 62952 -81210
rect 62706 -82361 62774 -82360
rect 62544 -82374 62600 -82364
rect 62720 -82370 62774 -82361
rect 62894 -81230 62898 -81220
rect 62950 -82368 62952 -82366
rect 62894 -82376 62952 -82368
rect 63056 -81218 63134 -81208
rect 63256 -81214 63310 -81204
rect 63056 -82364 63080 -81218
rect 63056 -82374 63134 -82364
rect 63254 -81228 63256 -81218
rect 62350 -82387 62404 -82376
rect 62894 -82378 62950 -82376
rect 63056 -82387 63110 -82374
rect 63254 -82376 63310 -82366
rect 63414 -81208 63468 -80744
rect 63622 -81206 63656 -81194
rect 63772 -81206 63826 -80744
rect 63978 -81204 64012 -81194
rect 64124 -81202 64178 -80744
rect 64468 -80886 66630 -80744
rect 63414 -81218 63486 -81208
rect 63414 -82364 63432 -81218
rect 63414 -82371 63486 -82364
rect 63432 -82374 63486 -82371
rect 63612 -81216 63666 -81206
rect 63772 -81216 63844 -81206
rect 63968 -81214 64022 -81204
rect 63666 -81230 63670 -81220
rect 63612 -82368 63614 -82362
rect 63612 -82372 63670 -82368
rect 63772 -82362 63790 -81216
rect 63772 -82371 63844 -82362
rect 63790 -82372 63844 -82371
rect 63966 -81224 63968 -81214
rect 63966 -82372 64022 -82362
rect 64124 -81212 64200 -81202
rect 64334 -81206 64368 -81196
rect 64124 -82358 64146 -81212
rect 64322 -81214 64376 -81206
rect 64124 -82368 64200 -82358
rect 64320 -81216 64376 -81214
rect 64320 -81224 64322 -81216
rect 63614 -82378 63670 -82372
rect 64124 -82383 64178 -82368
rect 64320 -82372 64376 -82362
rect 59568 -82442 59674 -82438
rect 62240 -82442 62346 -82438
rect 54804 -82448 64360 -82442
rect 54804 -82452 59568 -82448
rect 54804 -82608 56364 -82452
rect 56470 -82454 57086 -82452
rect 56470 -82458 56728 -82454
rect 56470 -82608 56546 -82458
rect 54804 -82614 56546 -82608
rect 56652 -82610 56728 -82458
rect 56834 -82610 56908 -82454
rect 57014 -82608 57086 -82454
rect 57192 -82608 57262 -82452
rect 57368 -82454 59390 -82452
rect 57368 -82608 57446 -82454
rect 57014 -82610 57446 -82608
rect 57552 -82610 57620 -82454
rect 57726 -82610 57794 -82454
rect 57900 -82458 58150 -82454
rect 57900 -82610 57976 -82458
rect 56652 -82614 57976 -82610
rect 58082 -82610 58150 -82458
rect 58256 -82610 58328 -82454
rect 58434 -82610 58508 -82454
rect 58614 -82610 58678 -82454
rect 58784 -82610 58858 -82454
rect 58964 -82610 59042 -82454
rect 59148 -82610 59216 -82454
rect 59322 -82608 59390 -82454
rect 59496 -82604 59568 -82452
rect 59674 -82454 62240 -82448
rect 59674 -82458 59926 -82454
rect 59674 -82604 59750 -82458
rect 59496 -82608 59750 -82604
rect 59322 -82610 59750 -82608
rect 58082 -82614 59750 -82610
rect 59856 -82610 59926 -82458
rect 60032 -82610 60106 -82454
rect 60212 -82610 60278 -82454
rect 60384 -82458 60636 -82454
rect 60384 -82610 60462 -82458
rect 59856 -82614 60462 -82610
rect 60568 -82610 60636 -82458
rect 60742 -82458 61168 -82454
rect 60742 -82610 60816 -82458
rect 60568 -82614 60816 -82610
rect 60922 -82614 60992 -82458
rect 61098 -82610 61168 -82458
rect 61274 -82458 61528 -82454
rect 61274 -82610 61348 -82458
rect 61098 -82614 61348 -82610
rect 61454 -82610 61528 -82458
rect 61634 -82462 61886 -82454
rect 61634 -82610 61706 -82462
rect 61454 -82614 61706 -82610
rect 54804 -82618 61706 -82614
rect 61812 -82610 61886 -82462
rect 61992 -82458 62240 -82454
rect 61992 -82610 62062 -82458
rect 61812 -82614 62062 -82610
rect 62168 -82604 62240 -82458
rect 62346 -82452 64360 -82448
rect 62346 -82454 63848 -82452
rect 62346 -82604 62418 -82454
rect 62168 -82610 62418 -82604
rect 62524 -82610 62596 -82454
rect 62702 -82458 63130 -82454
rect 62702 -82610 62776 -82458
rect 62168 -82614 62776 -82610
rect 62882 -82614 62956 -82458
rect 63062 -82610 63130 -82458
rect 63236 -82458 63848 -82454
rect 63236 -82610 63314 -82458
rect 63062 -82614 63314 -82610
rect 63420 -82614 63482 -82458
rect 63588 -82464 63848 -82458
rect 63588 -82614 63660 -82464
rect 61812 -82618 63660 -82614
rect 54804 -82620 63660 -82618
rect 63766 -82608 63848 -82464
rect 63954 -82454 64200 -82452
rect 63954 -82608 64020 -82454
rect 63766 -82610 64020 -82608
rect 64126 -82608 64200 -82454
rect 64306 -82608 64360 -82452
rect 64126 -82610 64360 -82608
rect 63766 -82620 64360 -82610
rect 54804 -82622 64360 -82620
rect 54810 -84294 54957 -82622
rect 56546 -82624 56652 -82622
rect 57976 -82624 58082 -82622
rect 59750 -82624 59856 -82622
rect 60462 -82624 60568 -82622
rect 60816 -82624 60922 -82622
rect 60992 -82624 61098 -82622
rect 61348 -82624 61454 -82622
rect 61706 -82628 61812 -82622
rect 62062 -82624 62168 -82622
rect 62776 -82624 62882 -82622
rect 62956 -82624 63062 -82622
rect 63314 -82624 63420 -82622
rect 63482 -82624 63588 -82622
rect 63660 -82630 63766 -82622
rect 56486 -82664 56520 -82656
rect 56842 -82664 56876 -82654
rect 56298 -82676 56352 -82666
rect 56474 -82670 56528 -82664
rect 56290 -83822 56298 -82683
rect 56290 -83832 56352 -83822
rect 56472 -82674 56528 -82670
rect 56472 -82680 56474 -82674
rect 56652 -82678 56706 -82668
rect 56472 -83820 56474 -83818
rect 56472 -83828 56528 -83820
rect 56474 -83830 56528 -83828
rect 56644 -83824 56652 -82689
rect 56486 -83832 56520 -83830
rect 53796 -84634 54958 -84294
rect 56290 -84314 56344 -83832
rect 56644 -83834 56706 -83824
rect 56836 -82674 56892 -82664
rect 56890 -83820 56892 -83812
rect 56836 -83822 56892 -83820
rect 57010 -82682 57064 -82672
rect 57198 -82676 57232 -82654
rect 57554 -82668 57588 -82654
rect 57542 -82670 57596 -82668
rect 56836 -83830 56890 -83822
rect 57180 -82686 57240 -82676
rect 57064 -83828 57066 -82699
rect 56644 -84314 56698 -83834
rect 57010 -83838 57066 -83828
rect 57366 -82682 57420 -82672
rect 57180 -83832 57186 -83824
rect 57180 -83834 57240 -83832
rect 57012 -84314 57066 -83838
rect 57186 -83842 57240 -83834
rect 57358 -83828 57366 -82689
rect 57540 -82678 57596 -82670
rect 57540 -82680 57542 -82678
rect 57724 -82678 57778 -82668
rect 57908 -82672 57942 -82656
rect 57540 -83824 57542 -83818
rect 57540 -83828 57596 -83824
rect 57358 -83838 57420 -83828
rect 57542 -83834 57596 -83828
rect 57716 -83824 57724 -82683
rect 57716 -83834 57778 -83824
rect 57900 -82676 57954 -82672
rect 57900 -82682 57956 -82676
rect 57954 -82686 57956 -82682
rect 58078 -82682 58132 -82672
rect 58266 -82676 58300 -82654
rect 58622 -82668 58656 -82654
rect 58978 -82668 59012 -82656
rect 59334 -82668 59368 -82654
rect 58260 -82678 58314 -82676
rect 57954 -83828 57956 -83824
rect 57900 -83834 57956 -83828
rect 58070 -83828 58078 -82683
rect 57358 -84314 57412 -83838
rect 57716 -84314 57770 -83834
rect 57900 -83838 57954 -83834
rect 58070 -83838 58132 -83828
rect 58258 -82686 58314 -82678
rect 58258 -82688 58260 -82686
rect 58258 -83832 58260 -83826
rect 58258 -83836 58314 -83832
rect 58070 -84314 58124 -83838
rect 58260 -83842 58314 -83836
rect 58434 -82682 58488 -82672
rect 58612 -82678 58668 -82668
rect 58612 -83826 58614 -83816
rect 58434 -84314 58488 -83828
rect 58614 -83836 58668 -83826
rect 58790 -82680 58844 -82670
rect 58970 -82672 59024 -82668
rect 58964 -82678 59024 -82672
rect 58964 -82682 58970 -82678
rect 58844 -83826 58846 -82683
rect 58790 -83836 58846 -83826
rect 59150 -82678 59204 -82668
rect 58964 -83824 58970 -83820
rect 58964 -83830 59024 -83824
rect 58970 -83834 59024 -83830
rect 59148 -83824 59150 -82683
rect 59148 -83834 59204 -83824
rect 59326 -82678 59382 -82668
rect 59506 -82673 59560 -82664
rect 59690 -82668 59724 -82654
rect 59682 -82672 59736 -82668
rect 60046 -82672 60080 -82656
rect 59326 -83824 59328 -83816
rect 59326 -83826 59382 -83824
rect 59328 -83834 59382 -83826
rect 59494 -82674 59560 -82673
rect 59494 -83820 59506 -82674
rect 59494 -83830 59560 -83820
rect 59678 -82678 59736 -82672
rect 59860 -82673 59914 -82672
rect 59678 -82682 59682 -82678
rect 59678 -83824 59682 -83820
rect 59678 -83830 59736 -83824
rect 58792 -84314 58846 -83836
rect 59148 -84314 59202 -83834
rect 59494 -84314 59548 -83830
rect 59682 -83834 59736 -83830
rect 59856 -82682 59914 -82673
rect 60038 -82680 60092 -82672
rect 59856 -83828 59860 -82682
rect 59856 -83838 59914 -83828
rect 60036 -82682 60092 -82680
rect 60036 -82690 60038 -82682
rect 60036 -83838 60092 -83828
rect 60212 -82682 60266 -82672
rect 60402 -82676 60436 -82658
rect 60758 -82668 60792 -82658
rect 60752 -82674 60806 -82668
rect 61114 -82672 61148 -82658
rect 61470 -82670 61504 -82658
rect 61462 -82672 61516 -82670
rect 60390 -82678 60444 -82676
rect 60386 -82686 60444 -82678
rect 60386 -82688 60390 -82686
rect 60266 -83828 60268 -82699
rect 60212 -83838 60268 -83828
rect 60572 -82686 60626 -82676
rect 60386 -83832 60390 -83826
rect 60386 -83836 60444 -83832
rect 59856 -84314 59910 -83838
rect 60214 -84314 60268 -83838
rect 60390 -83842 60444 -83836
rect 60560 -83832 60572 -82699
rect 60748 -82678 60806 -82674
rect 60748 -82684 60752 -82678
rect 60928 -82682 60982 -82672
rect 61106 -82678 61160 -82672
rect 60748 -83824 60752 -83822
rect 60748 -83832 60806 -83824
rect 60560 -83842 60626 -83832
rect 60752 -83834 60806 -83832
rect 60924 -83828 60928 -82721
rect 60924 -83838 60982 -83828
rect 61102 -82682 61160 -82678
rect 61102 -82688 61106 -82682
rect 61282 -82683 61336 -82676
rect 61102 -83828 61106 -83826
rect 61102 -83836 61160 -83828
rect 61106 -83838 61160 -83836
rect 61274 -82686 61336 -82683
rect 61274 -83832 61282 -82686
rect 61460 -82680 61516 -82672
rect 61460 -82682 61462 -82680
rect 61640 -82678 61694 -82668
rect 61826 -82672 61860 -82660
rect 62182 -82672 62216 -82662
rect 62538 -82670 62572 -82658
rect 61812 -82678 61866 -82672
rect 61460 -83826 61462 -83820
rect 61460 -83830 61516 -83826
rect 60560 -84314 60614 -83842
rect 60924 -84314 60978 -83838
rect 61274 -83842 61336 -83832
rect 61462 -83836 61516 -83830
rect 61632 -83824 61640 -82699
rect 61632 -83834 61694 -83824
rect 61810 -82682 61866 -82678
rect 61810 -82688 61812 -82682
rect 61810 -83828 61812 -83826
rect 61274 -84314 61328 -83842
rect 61632 -84314 61686 -83834
rect 61810 -83836 61866 -83828
rect 61812 -83838 61866 -83836
rect 61992 -82682 62046 -82672
rect 61992 -84314 62046 -83828
rect 62172 -82682 62226 -82672
rect 62352 -82682 62406 -82672
rect 62530 -82678 62584 -82670
rect 62226 -82692 62228 -82682
rect 62172 -83840 62228 -83830
rect 62338 -83828 62352 -82699
rect 62338 -83838 62406 -83828
rect 62528 -82680 62584 -82678
rect 62528 -82688 62530 -82680
rect 62528 -83836 62584 -83826
rect 62704 -82676 62758 -82666
rect 62894 -82672 62928 -82656
rect 63250 -82666 63284 -82656
rect 62882 -82682 62936 -82672
rect 62338 -84314 62392 -83838
rect 62704 -84314 62758 -83822
rect 62878 -82692 62882 -82682
rect 63064 -82680 63118 -82670
rect 63240 -82676 63294 -82666
rect 63606 -82668 63640 -82656
rect 63962 -82666 63996 -82656
rect 62934 -83830 62936 -83828
rect 62878 -83838 62936 -83830
rect 63060 -83826 63064 -82689
rect 63060 -83836 63118 -83826
rect 63238 -82690 63240 -82680
rect 63416 -82680 63470 -82670
rect 62878 -83840 62934 -83838
rect 63060 -84314 63114 -83836
rect 63238 -83838 63294 -83828
rect 63410 -83826 63416 -82699
rect 63410 -83836 63470 -83826
rect 63596 -82678 63650 -82668
rect 63774 -82678 63828 -82668
rect 63952 -82676 64006 -82666
rect 63650 -82692 63654 -82682
rect 63596 -83830 63598 -83824
rect 63596 -83834 63654 -83830
rect 63410 -84314 63464 -83836
rect 63598 -83840 63654 -83834
rect 63768 -83824 63774 -82689
rect 63768 -83834 63828 -83824
rect 63950 -82686 63952 -82676
rect 64130 -82674 64184 -82664
rect 64318 -82668 64352 -82658
rect 63950 -83834 64006 -83824
rect 64128 -83820 64130 -82683
rect 64306 -82676 64360 -82668
rect 64128 -83830 64184 -83820
rect 64304 -82678 64360 -82676
rect 64304 -82686 64306 -82678
rect 63768 -84314 63822 -83834
rect 64128 -84314 64182 -83830
rect 64304 -83834 64360 -83824
rect 64471 -83986 66630 -80886
rect 64468 -84314 66630 -83986
rect 56177 -84588 66630 -84314
rect 54810 -86258 54957 -84634
rect 56302 -85024 56356 -84588
rect 56474 -85022 56508 -85014
rect 56286 -85034 56356 -85024
rect 56462 -85028 56516 -85022
rect 56656 -85026 56710 -84588
rect 56830 -85022 56864 -85012
rect 56340 -86180 56356 -85034
rect 56286 -86190 56356 -86180
rect 56460 -85032 56516 -85028
rect 56460 -85038 56462 -85032
rect 56460 -86178 56462 -86176
rect 56460 -86186 56516 -86178
rect 56462 -86188 56516 -86186
rect 56640 -85036 56710 -85026
rect 56694 -86182 56710 -85036
rect 56474 -86190 56508 -86188
rect 56302 -86205 56356 -86190
rect 56640 -86192 56710 -86182
rect 56824 -85032 56880 -85022
rect 57012 -85030 57066 -84588
rect 56878 -86178 56880 -86170
rect 56824 -86180 56880 -86178
rect 56998 -85040 57066 -85030
rect 57186 -85034 57220 -85012
rect 57370 -85030 57424 -84588
rect 57542 -85026 57576 -85012
rect 57720 -85026 57774 -84588
rect 57530 -85028 57584 -85026
rect 56824 -86188 56878 -86180
rect 57052 -86186 57066 -85040
rect 56656 -86193 56710 -86192
rect 56998 -86193 57066 -86186
rect 57168 -85044 57228 -85034
rect 57168 -86190 57174 -86182
rect 57168 -86192 57228 -86190
rect 56998 -86196 57052 -86193
rect 57174 -86200 57228 -86192
rect 57354 -85040 57424 -85030
rect 57408 -86186 57424 -85040
rect 57528 -85036 57584 -85028
rect 57528 -85038 57530 -85036
rect 57528 -86182 57530 -86176
rect 57528 -86186 57584 -86182
rect 57354 -86196 57424 -86186
rect 57530 -86192 57584 -86186
rect 57712 -85036 57774 -85026
rect 57896 -85030 57930 -85014
rect 58084 -85030 58138 -84588
rect 57766 -86182 57774 -85036
rect 57712 -86192 57774 -86182
rect 57370 -86209 57424 -86196
rect 57720 -86209 57774 -86192
rect 57888 -85034 57942 -85030
rect 57888 -85040 57944 -85034
rect 57942 -85044 57944 -85040
rect 57942 -86186 57944 -86182
rect 57888 -86192 57944 -86186
rect 58066 -85040 58138 -85030
rect 58254 -85034 58288 -85012
rect 58434 -85030 58488 -84588
rect 58610 -85026 58644 -85012
rect 58248 -85036 58302 -85034
rect 58120 -86186 58138 -85040
rect 57888 -86196 57942 -86192
rect 58066 -86196 58138 -86186
rect 58246 -85044 58302 -85036
rect 58246 -85046 58248 -85044
rect 58246 -86190 58248 -86184
rect 58246 -86194 58302 -86190
rect 58084 -86221 58138 -86196
rect 58248 -86200 58302 -86194
rect 58422 -85040 58488 -85030
rect 58476 -86186 58488 -85040
rect 58600 -85036 58656 -85026
rect 58792 -85028 58846 -84588
rect 58966 -85026 59000 -85014
rect 59148 -85026 59202 -84588
rect 59322 -85026 59356 -85012
rect 59498 -85022 59552 -84588
rect 58600 -86184 58602 -86174
rect 58422 -86193 58488 -86186
rect 58422 -86196 58476 -86193
rect 58602 -86194 58656 -86184
rect 58778 -85038 58846 -85028
rect 58958 -85030 59012 -85026
rect 58832 -86177 58846 -85038
rect 58952 -85036 59012 -85030
rect 58952 -85040 58958 -85036
rect 58778 -86194 58832 -86184
rect 58952 -86182 58958 -86178
rect 58952 -86188 59012 -86182
rect 58958 -86192 59012 -86188
rect 59138 -85036 59202 -85026
rect 59192 -86182 59202 -85036
rect 59138 -86183 59202 -86182
rect 59314 -85036 59370 -85026
rect 59314 -86182 59316 -86174
rect 59138 -86192 59192 -86183
rect 59314 -86184 59370 -86182
rect 59316 -86192 59370 -86184
rect 59494 -85032 59552 -85022
rect 59678 -85026 59712 -85012
rect 59670 -85030 59724 -85026
rect 59864 -85030 59918 -84588
rect 60034 -85030 60068 -85014
rect 60210 -85030 60264 -84588
rect 59548 -86167 59552 -85032
rect 59666 -85036 59724 -85030
rect 59666 -85040 59670 -85036
rect 59494 -86188 59548 -86178
rect 59666 -86182 59670 -86178
rect 59666 -86188 59724 -86182
rect 59670 -86192 59724 -86188
rect 59848 -85040 59918 -85030
rect 60026 -85038 60080 -85030
rect 59902 -86186 59918 -85040
rect 59848 -86196 59918 -86186
rect 60024 -85040 60080 -85038
rect 60024 -85048 60026 -85040
rect 60024 -86196 60080 -86186
rect 60200 -85040 60264 -85030
rect 60390 -85034 60424 -85016
rect 60570 -85034 60624 -84588
rect 60746 -85026 60780 -85016
rect 60740 -85032 60794 -85026
rect 60928 -85030 60982 -84588
rect 61102 -85030 61136 -85016
rect 60378 -85036 60432 -85034
rect 60254 -86186 60264 -85040
rect 60200 -86196 60264 -86186
rect 60374 -85044 60432 -85036
rect 60374 -85046 60378 -85044
rect 60374 -86190 60378 -86184
rect 60374 -86194 60432 -86190
rect 59864 -86205 59918 -86196
rect 60210 -86221 60264 -86196
rect 60378 -86200 60432 -86194
rect 60560 -85044 60624 -85034
rect 60614 -86183 60624 -85044
rect 60736 -85036 60794 -85032
rect 60736 -85042 60740 -85036
rect 60736 -86182 60740 -86180
rect 60736 -86190 60794 -86182
rect 60560 -86200 60614 -86190
rect 60740 -86192 60794 -86190
rect 60916 -85040 60982 -85030
rect 61094 -85036 61148 -85030
rect 61282 -85034 61336 -84588
rect 61458 -85028 61492 -85016
rect 61638 -85026 61692 -84588
rect 61450 -85030 61504 -85028
rect 60970 -86186 60982 -85040
rect 60916 -86193 60982 -86186
rect 61090 -85040 61148 -85036
rect 61090 -85046 61094 -85040
rect 61090 -86186 61094 -86184
rect 60916 -86196 60970 -86193
rect 61090 -86194 61148 -86186
rect 61094 -86196 61148 -86194
rect 61270 -85044 61336 -85034
rect 61324 -86190 61336 -85044
rect 61448 -85038 61504 -85030
rect 61448 -85040 61450 -85038
rect 61448 -86184 61450 -86178
rect 61448 -86188 61504 -86184
rect 61270 -86200 61336 -86190
rect 61450 -86194 61504 -86188
rect 61628 -85036 61692 -85026
rect 61814 -85030 61848 -85018
rect 61996 -85030 62050 -84588
rect 62170 -85030 62204 -85020
rect 62354 -85030 62408 -84588
rect 62526 -85028 62560 -85016
rect 62710 -85024 62764 -84588
rect 61800 -85036 61854 -85030
rect 61682 -86182 61692 -85036
rect 61628 -86183 61692 -86182
rect 61798 -85040 61854 -85036
rect 61798 -85046 61800 -85040
rect 61628 -86192 61682 -86183
rect 61798 -86186 61800 -86184
rect 61798 -86194 61854 -86186
rect 61800 -86196 61854 -86194
rect 61980 -85040 62050 -85030
rect 62034 -86186 62050 -85040
rect 61980 -86196 62050 -86186
rect 61282 -86209 61336 -86200
rect 61996 -86209 62050 -86196
rect 62160 -85040 62214 -85030
rect 62340 -85040 62408 -85030
rect 62518 -85036 62572 -85028
rect 62214 -85050 62216 -85040
rect 62160 -86198 62216 -86188
rect 62394 -86186 62408 -85040
rect 62340 -86196 62408 -86186
rect 62516 -85038 62572 -85036
rect 62516 -85046 62518 -85038
rect 62516 -86194 62572 -86184
rect 62692 -85034 62764 -85024
rect 62882 -85030 62916 -85014
rect 63060 -85028 63114 -84588
rect 63238 -85024 63272 -85014
rect 62746 -86180 62764 -85034
rect 62870 -85040 62924 -85030
rect 62692 -86183 62764 -86180
rect 62866 -85050 62870 -85040
rect 62692 -86190 62746 -86183
rect 62922 -86188 62924 -86186
rect 62354 -86209 62408 -86196
rect 62866 -86196 62924 -86188
rect 63052 -85038 63114 -85028
rect 63228 -85034 63282 -85024
rect 63418 -85028 63472 -84588
rect 63594 -85026 63628 -85014
rect 63776 -85026 63830 -84588
rect 63950 -85024 63984 -85014
rect 64128 -85022 64182 -84588
rect 63106 -86184 63114 -85038
rect 63052 -86193 63114 -86184
rect 63226 -85048 63228 -85038
rect 63052 -86194 63106 -86193
rect 63226 -86196 63282 -86186
rect 63404 -85038 63472 -85028
rect 63458 -86184 63472 -85038
rect 63404 -86194 63472 -86184
rect 63584 -85036 63638 -85026
rect 63762 -85036 63830 -85026
rect 63940 -85034 63994 -85024
rect 63638 -85050 63642 -85040
rect 63584 -86188 63586 -86182
rect 63584 -86192 63642 -86188
rect 63816 -86182 63830 -85036
rect 63762 -86192 63830 -86182
rect 63938 -85044 63940 -85034
rect 63938 -86192 63994 -86182
rect 64118 -85032 64182 -85022
rect 64306 -85026 64340 -85016
rect 64172 -86177 64182 -85032
rect 64294 -85034 64348 -85026
rect 64292 -85036 64348 -85034
rect 64292 -85044 64294 -85036
rect 64118 -86188 64172 -86178
rect 64292 -86192 64348 -86182
rect 62866 -86198 62922 -86196
rect 63418 -86227 63472 -86194
rect 63586 -86198 63642 -86192
rect 63776 -86209 63830 -86192
rect 54810 -86268 64346 -86258
rect 54810 -86272 59540 -86268
rect 54810 -86428 56336 -86272
rect 56442 -86274 57058 -86272
rect 56442 -86278 56700 -86274
rect 56442 -86428 56518 -86278
rect 54810 -86434 56518 -86428
rect 56624 -86430 56700 -86278
rect 56806 -86430 56880 -86274
rect 56986 -86428 57058 -86274
rect 57164 -86428 57234 -86272
rect 57340 -86274 59362 -86272
rect 57340 -86428 57418 -86274
rect 56986 -86430 57418 -86428
rect 57524 -86430 57592 -86274
rect 57698 -86430 57766 -86274
rect 57872 -86278 58122 -86274
rect 57872 -86430 57948 -86278
rect 56624 -86434 57948 -86430
rect 58054 -86430 58122 -86278
rect 58228 -86430 58300 -86274
rect 58406 -86430 58480 -86274
rect 58586 -86430 58650 -86274
rect 58756 -86430 58830 -86274
rect 58936 -86430 59014 -86274
rect 59120 -86430 59188 -86274
rect 59294 -86428 59362 -86274
rect 59468 -86424 59540 -86272
rect 59646 -86274 62212 -86268
rect 59646 -86278 59898 -86274
rect 59646 -86424 59722 -86278
rect 59468 -86428 59722 -86424
rect 59294 -86430 59722 -86428
rect 58054 -86434 59722 -86430
rect 59828 -86430 59898 -86278
rect 60004 -86430 60078 -86274
rect 60184 -86430 60250 -86274
rect 60356 -86278 60608 -86274
rect 60356 -86430 60434 -86278
rect 59828 -86434 60434 -86430
rect 60540 -86430 60608 -86278
rect 60714 -86278 61140 -86274
rect 60714 -86430 60788 -86278
rect 60540 -86434 60788 -86430
rect 60894 -86434 60964 -86278
rect 61070 -86430 61140 -86278
rect 61246 -86278 61500 -86274
rect 61246 -86430 61320 -86278
rect 61070 -86434 61320 -86430
rect 61426 -86430 61500 -86278
rect 61606 -86282 61858 -86274
rect 61606 -86430 61678 -86282
rect 61426 -86434 61678 -86430
rect 54810 -86438 61678 -86434
rect 61784 -86430 61858 -86282
rect 61964 -86278 62212 -86274
rect 61964 -86430 62034 -86278
rect 61784 -86434 62034 -86430
rect 62140 -86424 62212 -86278
rect 62318 -86272 64346 -86268
rect 62318 -86274 63820 -86272
rect 62318 -86424 62390 -86274
rect 62140 -86430 62390 -86424
rect 62496 -86430 62568 -86274
rect 62674 -86278 63102 -86274
rect 62674 -86430 62748 -86278
rect 62140 -86434 62748 -86430
rect 62854 -86434 62928 -86278
rect 63034 -86430 63102 -86278
rect 63208 -86278 63820 -86274
rect 63208 -86430 63286 -86278
rect 63034 -86434 63286 -86430
rect 63392 -86434 63454 -86278
rect 63560 -86284 63820 -86278
rect 63560 -86434 63632 -86284
rect 61784 -86438 63632 -86434
rect 56518 -86444 56624 -86438
rect 56700 -86440 56806 -86438
rect 56880 -86440 56986 -86438
rect 57418 -86440 57524 -86438
rect 57592 -86440 57698 -86438
rect 57766 -86440 57872 -86438
rect 57948 -86444 58054 -86438
rect 58122 -86440 58228 -86438
rect 58300 -86440 58406 -86438
rect 58480 -86440 58586 -86438
rect 58650 -86440 58756 -86438
rect 58830 -86440 58936 -86438
rect 59014 -86440 59120 -86438
rect 59188 -86440 59294 -86438
rect 59722 -86444 59828 -86438
rect 59898 -86440 60004 -86438
rect 60078 -86440 60184 -86438
rect 60250 -86440 60356 -86438
rect 60434 -86444 60540 -86438
rect 60608 -86440 60714 -86438
rect 60788 -86444 60894 -86438
rect 60964 -86444 61070 -86438
rect 61140 -86440 61246 -86438
rect 61320 -86444 61426 -86438
rect 61500 -86440 61606 -86438
rect 61678 -86448 61784 -86438
rect 61858 -86440 61964 -86438
rect 62034 -86444 62140 -86438
rect 62390 -86440 62496 -86438
rect 62568 -86440 62674 -86438
rect 62748 -86444 62854 -86438
rect 62928 -86444 63034 -86438
rect 63102 -86440 63208 -86438
rect 63286 -86444 63392 -86438
rect 63454 -86444 63560 -86438
rect 63738 -86428 63820 -86284
rect 63926 -86274 64172 -86272
rect 63926 -86428 63992 -86274
rect 63738 -86430 63992 -86428
rect 64098 -86428 64172 -86274
rect 64278 -86428 64346 -86272
rect 64098 -86430 64346 -86428
rect 63738 -86438 64346 -86430
rect 64468 -86422 66630 -84588
rect 63992 -86440 64098 -86438
rect 63632 -86450 63738 -86440
rect 56458 -86484 56492 -86476
rect 56814 -86484 56848 -86474
rect 56270 -86496 56324 -86486
rect 56446 -86490 56500 -86484
rect 56444 -86494 56500 -86490
rect 56444 -86500 56446 -86494
rect 56324 -87642 56348 -86505
rect 56270 -87652 56348 -87642
rect 56444 -87640 56446 -87638
rect 56444 -87648 56500 -87640
rect 56446 -87650 56500 -87648
rect 56624 -86498 56678 -86488
rect 56808 -86494 56864 -86484
rect 56678 -87644 56702 -86511
rect 56458 -87652 56492 -87650
rect 55742 -87954 56040 -87944
rect 56294 -88024 56348 -87652
rect 56624 -87654 56702 -87644
rect 56862 -87640 56864 -87632
rect 56808 -87642 56864 -87640
rect 56982 -86495 57036 -86492
rect 56982 -86502 57070 -86495
rect 57170 -86496 57204 -86474
rect 57526 -86488 57560 -86474
rect 57514 -86490 57568 -86488
rect 57338 -86495 57392 -86492
rect 56808 -87650 56862 -87642
rect 57036 -87648 57070 -86502
rect 56648 -88024 56702 -87654
rect 56982 -87658 57070 -87648
rect 57152 -86506 57212 -86496
rect 57152 -87652 57158 -87644
rect 57152 -87654 57212 -87652
rect 57016 -88024 57070 -87658
rect 57158 -87662 57212 -87654
rect 57338 -86502 57416 -86495
rect 57392 -87648 57416 -86502
rect 57512 -86498 57568 -86490
rect 57512 -86500 57514 -86498
rect 57512 -87644 57514 -87638
rect 57512 -87648 57568 -87644
rect 57338 -87658 57416 -87648
rect 57514 -87654 57568 -87648
rect 57696 -86495 57750 -86488
rect 57880 -86492 57914 -86476
rect 57696 -86498 57774 -86495
rect 57750 -87644 57774 -86498
rect 57696 -87654 57774 -87644
rect 57362 -88024 57416 -87658
rect 57720 -88024 57774 -87654
rect 57872 -86496 57926 -86492
rect 58050 -86495 58104 -86492
rect 57872 -86502 57928 -86496
rect 57926 -86506 57928 -86502
rect 57926 -87648 57928 -87644
rect 57872 -87654 57928 -87648
rect 58050 -86502 58128 -86495
rect 58238 -86496 58272 -86474
rect 58594 -86488 58628 -86474
rect 58950 -86488 58984 -86476
rect 59306 -86488 59340 -86474
rect 58232 -86498 58286 -86496
rect 58104 -87648 58128 -86502
rect 57872 -87658 57926 -87654
rect 58050 -87658 58128 -87648
rect 58230 -86506 58286 -86498
rect 58230 -86508 58232 -86506
rect 58230 -87652 58232 -87646
rect 58230 -87656 58286 -87652
rect 58074 -88024 58128 -87658
rect 58232 -87662 58286 -87656
rect 58406 -86502 58460 -86492
rect 58584 -86498 58640 -86488
rect 58460 -87648 58492 -86511
rect 58584 -87646 58586 -87636
rect 58406 -87658 58492 -87648
rect 58586 -87656 58640 -87646
rect 58762 -86500 58816 -86490
rect 58942 -86492 58996 -86488
rect 58936 -86498 58996 -86492
rect 58936 -86502 58942 -86498
rect 58816 -87646 58850 -86505
rect 58762 -87656 58850 -87646
rect 58936 -87644 58942 -87640
rect 58936 -87650 58996 -87644
rect 58942 -87654 58996 -87650
rect 59122 -86498 59176 -86488
rect 59298 -86498 59354 -86488
rect 59176 -87644 59206 -86505
rect 59122 -87654 59206 -87644
rect 59298 -87644 59300 -87636
rect 59298 -87646 59354 -87644
rect 59300 -87654 59354 -87646
rect 59478 -86494 59532 -86484
rect 59662 -86488 59696 -86474
rect 59654 -86492 59708 -86488
rect 60018 -86492 60052 -86476
rect 59650 -86498 59708 -86492
rect 59650 -86502 59654 -86498
rect 59532 -87640 59552 -86511
rect 59478 -87650 59552 -87640
rect 59650 -87644 59654 -87640
rect 59650 -87650 59708 -87644
rect 58438 -88024 58492 -87658
rect 58796 -88024 58850 -87656
rect 59152 -88024 59206 -87654
rect 59498 -88024 59552 -87650
rect 59654 -87654 59708 -87650
rect 59832 -86502 59886 -86492
rect 60010 -86500 60064 -86492
rect 60008 -86502 60064 -86500
rect 60008 -86510 60010 -86502
rect 59886 -87648 59914 -86511
rect 59832 -87658 59914 -87648
rect 60008 -87658 60064 -87648
rect 60184 -86502 60238 -86492
rect 60374 -86496 60408 -86478
rect 60730 -86488 60764 -86478
rect 60724 -86494 60778 -86488
rect 61086 -86492 61120 -86478
rect 61442 -86490 61476 -86478
rect 61434 -86492 61488 -86490
rect 60362 -86498 60416 -86496
rect 60238 -87648 60272 -86505
rect 60184 -87658 60272 -87648
rect 60358 -86506 60416 -86498
rect 60358 -86508 60362 -86506
rect 60358 -87652 60362 -87646
rect 60358 -87656 60416 -87652
rect 59860 -88024 59914 -87658
rect 60218 -88024 60272 -87658
rect 60362 -87662 60416 -87656
rect 60544 -86505 60598 -86496
rect 60720 -86498 60778 -86494
rect 60720 -86504 60724 -86498
rect 60544 -86506 60618 -86505
rect 60598 -87652 60618 -86506
rect 60720 -87644 60724 -87642
rect 60720 -87652 60778 -87644
rect 60544 -87662 60618 -87652
rect 60724 -87654 60778 -87652
rect 60900 -86502 60954 -86492
rect 61078 -86498 61132 -86492
rect 61278 -86496 61332 -86495
rect 61074 -86502 61132 -86498
rect 60954 -87648 60982 -86505
rect 60900 -87658 60982 -87648
rect 61074 -86508 61078 -86502
rect 61074 -87648 61078 -87646
rect 61074 -87656 61132 -87648
rect 61078 -87658 61132 -87656
rect 61254 -86506 61332 -86496
rect 61308 -87652 61332 -86506
rect 61432 -86500 61488 -86492
rect 61432 -86502 61434 -86500
rect 61432 -87646 61434 -87640
rect 61432 -87650 61488 -87646
rect 60564 -88024 60618 -87662
rect 60928 -88024 60982 -87658
rect 61254 -87662 61332 -87652
rect 61434 -87656 61488 -87650
rect 61612 -86498 61666 -86488
rect 61798 -86492 61832 -86480
rect 62154 -86492 62188 -86482
rect 62510 -86490 62544 -86478
rect 61784 -86498 61838 -86492
rect 61782 -86502 61838 -86498
rect 61782 -86508 61784 -86502
rect 61666 -87644 61690 -86511
rect 61612 -87654 61690 -87644
rect 61278 -88024 61332 -87662
rect 61636 -88024 61690 -87654
rect 61782 -87648 61784 -87646
rect 61782 -87656 61838 -87648
rect 61784 -87658 61838 -87656
rect 61964 -86495 62018 -86492
rect 61964 -86502 62050 -86495
rect 62018 -87648 62050 -86502
rect 61964 -87658 62050 -87648
rect 61996 -88024 62050 -87658
rect 62144 -86502 62198 -86492
rect 62324 -86495 62378 -86492
rect 62324 -86502 62396 -86495
rect 62502 -86498 62556 -86490
rect 62198 -86512 62200 -86502
rect 62144 -87660 62200 -87650
rect 62378 -87648 62396 -86502
rect 62324 -87658 62396 -87648
rect 62500 -86500 62556 -86498
rect 62500 -86508 62502 -86500
rect 62500 -87656 62556 -87646
rect 62676 -86495 62730 -86486
rect 62866 -86492 62900 -86476
rect 63222 -86486 63256 -86476
rect 62676 -86496 62762 -86495
rect 62730 -87642 62762 -86496
rect 62854 -86502 62908 -86492
rect 62676 -87652 62762 -87642
rect 62342 -88024 62396 -87658
rect 62708 -88024 62762 -87652
rect 62850 -86512 62854 -86502
rect 62906 -87650 62908 -87648
rect 62850 -87658 62908 -87650
rect 63036 -86495 63090 -86490
rect 63036 -86500 63118 -86495
rect 63212 -86496 63266 -86486
rect 63414 -86490 63468 -86483
rect 63578 -86488 63612 -86476
rect 63934 -86486 63968 -86476
rect 63090 -87646 63118 -86500
rect 63036 -87656 63118 -87646
rect 62850 -87660 62906 -87658
rect 63064 -88024 63118 -87656
rect 63210 -86510 63212 -86500
rect 63210 -87658 63266 -87648
rect 63388 -86500 63468 -86490
rect 63442 -87646 63468 -86500
rect 63388 -87656 63468 -87646
rect 63568 -86498 63622 -86488
rect 63746 -86495 63800 -86488
rect 63746 -86498 63826 -86495
rect 63924 -86496 63978 -86486
rect 63622 -86512 63626 -86502
rect 63568 -87650 63570 -87644
rect 63568 -87654 63626 -87650
rect 63800 -87644 63826 -86498
rect 63746 -87654 63826 -87644
rect 63922 -86506 63924 -86496
rect 63922 -87654 63978 -87644
rect 64102 -86494 64156 -86484
rect 64290 -86488 64324 -86478
rect 64156 -87640 64186 -86495
rect 64278 -86496 64332 -86488
rect 64102 -87650 64186 -87640
rect 63414 -88024 63468 -87656
rect 63570 -87660 63626 -87654
rect 63772 -88024 63826 -87654
rect 64132 -88024 64186 -87650
rect 64276 -86498 64332 -86496
rect 64276 -86506 64278 -86498
rect 64276 -87654 64332 -87644
rect 64468 -88024 65484 -86422
rect 56040 -88298 65484 -88024
rect 64964 -88304 65484 -88298
rect 65906 -87278 66524 -87042
rect 65906 -87398 66526 -87278
rect 65906 -87842 66042 -87398
rect 66108 -87442 67286 -87440
rect 66108 -87534 67842 -87442
rect 66108 -87574 67286 -87534
rect 66154 -87606 66188 -87574
rect 66510 -87602 66544 -87574
rect 66140 -87616 66196 -87606
rect 66318 -87614 66374 -87604
rect 66140 -87800 66196 -87790
rect 66316 -87634 66318 -87624
rect 66316 -87798 66374 -87788
rect 66498 -87612 66554 -87602
rect 66866 -87604 66900 -87574
rect 67222 -87602 67256 -87574
rect 66676 -87614 66732 -87604
rect 66498 -87796 66554 -87786
rect 66674 -87634 66676 -87624
rect 66674 -87798 66732 -87788
rect 66848 -87614 66904 -87604
rect 67030 -87612 67086 -87602
rect 66848 -87798 66904 -87788
rect 67028 -87632 67030 -87622
rect 67028 -87796 67086 -87786
rect 67208 -87612 67264 -87602
rect 67208 -87796 67264 -87786
rect 66212 -87838 66316 -87828
rect 65906 -87988 66212 -87842
rect 55742 -88364 56040 -88354
rect 54816 -89040 65498 -88610
rect 65906 -88684 66042 -87988
rect 66392 -87838 66496 -87828
rect 66316 -87988 66392 -87842
rect 66212 -88000 66316 -87990
rect 66570 -87838 66674 -87828
rect 66496 -87988 66570 -87842
rect 66392 -88000 66496 -87990
rect 66746 -87838 66850 -87828
rect 66674 -87988 66746 -87842
rect 66570 -88000 66674 -87990
rect 66924 -87838 67028 -87828
rect 66850 -87988 66924 -87842
rect 66746 -88000 66850 -87990
rect 67100 -87838 67204 -87828
rect 67028 -87988 67100 -87842
rect 66924 -88000 67028 -87990
rect 67204 -87988 67276 -87842
rect 67100 -88000 67204 -87990
rect 66146 -88044 66202 -88034
rect 66326 -88040 66382 -88030
rect 66146 -88228 66202 -88218
rect 66324 -88060 66326 -88050
rect 66324 -88224 66382 -88214
rect 66506 -88042 66562 -88032
rect 66506 -88226 66562 -88216
rect 66684 -88042 66740 -88032
rect 66862 -88042 66918 -88032
rect 66740 -88070 66758 -88060
rect 66684 -88224 66702 -88216
rect 66684 -88226 66758 -88224
rect 67040 -88042 67096 -88032
rect 66862 -88226 66918 -88216
rect 67038 -88062 67040 -88052
rect 67038 -88226 67096 -88216
rect 67218 -88046 67274 -88036
rect 66154 -88314 66188 -88228
rect 66510 -88314 66544 -88226
rect 66702 -88234 66758 -88226
rect 66866 -88314 66900 -88226
rect 67218 -88230 67274 -88220
rect 67222 -88314 67256 -88230
rect 67554 -88314 67842 -87534
rect 80284 -87854 80318 -87850
rect 68274 -87862 68308 -87858
rect 66108 -88362 67842 -88314
rect 66154 -88442 66188 -88362
rect 66136 -88452 66192 -88442
rect 66320 -88446 66376 -88436
rect 66510 -88440 66544 -88362
rect 66866 -88436 66900 -88362
rect 66136 -88636 66192 -88626
rect 66318 -88466 66320 -88456
rect 66318 -88630 66376 -88620
rect 66500 -88450 66556 -88440
rect 66676 -88452 66732 -88442
rect 66332 -88632 66366 -88630
rect 66500 -88634 66556 -88624
rect 66674 -88472 66676 -88462
rect 66674 -88636 66732 -88626
rect 66854 -88446 66910 -88436
rect 67034 -88448 67090 -88438
rect 67222 -88442 67256 -88362
rect 66854 -88630 66910 -88620
rect 67032 -88468 67034 -88458
rect 66866 -88632 66900 -88630
rect 67032 -88632 67090 -88622
rect 67212 -88452 67268 -88442
rect 67212 -88636 67268 -88626
rect 66210 -88674 66314 -88664
rect 65906 -88826 66210 -88684
rect 66392 -88676 66496 -88666
rect 66314 -88826 66392 -88684
rect 65906 -88828 66392 -88826
rect 66564 -88678 66668 -88668
rect 66496 -88828 66564 -88684
rect 65906 -88830 66564 -88828
rect 66746 -88678 66850 -88668
rect 66668 -88830 66746 -88684
rect 66924 -88678 67028 -88668
rect 66850 -88830 66924 -88684
rect 67104 -88678 67208 -88668
rect 67028 -88830 67104 -88684
rect 67208 -88830 67294 -88684
rect 66210 -88836 66314 -88830
rect 66392 -88838 66496 -88830
rect 66564 -88840 66668 -88830
rect 66746 -88840 66850 -88830
rect 66924 -88840 67028 -88830
rect 67104 -88840 67208 -88830
rect 66140 -88874 66192 -88864
rect 54816 -89042 65318 -89040
rect 54816 -89050 64644 -89042
rect 54816 -90632 55860 -89050
rect 66140 -89073 66192 -89028
rect 66318 -88880 66374 -88870
rect 66318 -89044 66374 -89034
rect 66496 -88876 66548 -88866
rect 66496 -89040 66548 -89030
rect 66670 -88880 66726 -88870
rect 66510 -89073 66544 -89040
rect 66670 -89044 66726 -89034
rect 66852 -88882 66904 -88872
rect 66852 -89046 66904 -89036
rect 67032 -88880 67088 -88870
rect 67224 -88873 67276 -88872
rect 67032 -89044 67088 -89034
rect 67222 -88882 67276 -88873
rect 67222 -89036 67224 -88882
rect 67222 -89046 67276 -89036
rect 66107 -89074 66544 -89073
rect 66866 -89074 66900 -89046
rect 67222 -89074 67256 -89046
rect 67554 -89074 67842 -88362
rect 68260 -87872 68318 -87862
rect 68260 -89034 68318 -89024
rect 68440 -87868 68498 -87858
rect 68440 -89030 68498 -89020
rect 68628 -87868 68686 -87858
rect 68808 -87864 68842 -87858
rect 68986 -87862 69020 -87858
rect 68628 -89030 68686 -89020
rect 68802 -87874 68860 -87864
rect 68452 -89034 68486 -89030
rect 68630 -89034 68664 -89030
rect 68802 -89036 68860 -89026
rect 68978 -87872 69036 -87862
rect 69164 -87864 69198 -87858
rect 69342 -87864 69376 -87858
rect 69520 -87862 69554 -87858
rect 69698 -87862 69732 -87858
rect 68978 -89026 68980 -89024
rect 69032 -89026 69036 -89024
rect 68978 -89034 69036 -89026
rect 69160 -87874 69218 -87864
rect 69338 -87874 69396 -87864
rect 68980 -89036 69032 -89034
rect 69160 -89036 69218 -89026
rect 69336 -87890 69338 -87880
rect 69336 -89036 69396 -89026
rect 69512 -87872 69570 -87862
rect 69512 -89034 69570 -89024
rect 69692 -87872 69750 -87862
rect 69876 -87864 69910 -87858
rect 69692 -89034 69750 -89024
rect 69866 -87874 69924 -87864
rect 70054 -87868 70088 -87858
rect 69866 -89036 69924 -89026
rect 70048 -87878 70106 -87868
rect 70232 -87870 70266 -87858
rect 70410 -87862 70444 -87858
rect 70048 -89040 70106 -89030
rect 70222 -87880 70280 -87870
rect 70222 -89042 70280 -89032
rect 70400 -87872 70458 -87862
rect 70588 -87868 70622 -87858
rect 70766 -87868 70800 -87858
rect 70944 -87866 70978 -87858
rect 71122 -87866 71156 -87858
rect 70400 -89034 70458 -89024
rect 70582 -87878 70640 -87868
rect 70582 -89040 70640 -89030
rect 70756 -87878 70814 -87868
rect 70756 -89040 70814 -89030
rect 70936 -87876 70994 -87866
rect 71118 -87876 71176 -87866
rect 71300 -87872 71334 -87858
rect 71478 -87870 71512 -87858
rect 71656 -87870 71690 -87858
rect 71834 -87866 71868 -87858
rect 74170 -87860 74204 -87856
rect 70936 -89038 70994 -89028
rect 71114 -87892 71118 -87882
rect 71114 -89038 71176 -89028
rect 71292 -87882 71350 -87872
rect 71292 -89044 71350 -89034
rect 71472 -87880 71530 -87870
rect 71472 -89042 71530 -89032
rect 71646 -87880 71704 -87870
rect 71646 -89042 71704 -89032
rect 71824 -87876 71882 -87866
rect 71824 -89038 71882 -89028
rect 74156 -87870 74214 -87860
rect 74156 -89032 74214 -89022
rect 74336 -87866 74394 -87856
rect 74336 -89028 74394 -89018
rect 74524 -87866 74582 -87856
rect 74704 -87862 74738 -87856
rect 74882 -87860 74916 -87856
rect 74524 -89028 74582 -89018
rect 74698 -87872 74756 -87862
rect 74348 -89032 74382 -89028
rect 74526 -89032 74560 -89028
rect 74698 -89034 74756 -89024
rect 74874 -87870 74932 -87860
rect 75060 -87862 75094 -87856
rect 75238 -87862 75272 -87856
rect 75416 -87860 75450 -87856
rect 75594 -87860 75628 -87856
rect 74874 -89024 74876 -89022
rect 74928 -89024 74932 -89022
rect 74874 -89032 74932 -89024
rect 75056 -87872 75114 -87862
rect 75234 -87872 75292 -87862
rect 74876 -89034 74928 -89032
rect 75056 -89034 75114 -89024
rect 75232 -87888 75234 -87878
rect 75232 -89034 75292 -89024
rect 75408 -87870 75466 -87860
rect 75408 -89032 75466 -89022
rect 75588 -87870 75646 -87860
rect 75772 -87862 75806 -87856
rect 75588 -89032 75646 -89022
rect 75762 -87872 75820 -87862
rect 75950 -87866 75984 -87856
rect 75762 -89034 75820 -89024
rect 75944 -87876 76002 -87866
rect 76128 -87868 76162 -87856
rect 76306 -87860 76340 -87856
rect 75944 -89038 76002 -89028
rect 76118 -87878 76176 -87868
rect 76118 -89040 76176 -89030
rect 76296 -87870 76354 -87860
rect 76484 -87866 76518 -87856
rect 76662 -87866 76696 -87856
rect 76840 -87864 76874 -87856
rect 77018 -87864 77052 -87856
rect 76296 -89032 76354 -89022
rect 76478 -87876 76536 -87866
rect 76478 -89038 76536 -89028
rect 76652 -87876 76710 -87866
rect 76652 -89038 76710 -89028
rect 76832 -87874 76890 -87864
rect 77014 -87874 77072 -87864
rect 77196 -87870 77230 -87856
rect 77374 -87868 77408 -87856
rect 77552 -87868 77586 -87856
rect 77730 -87864 77764 -87856
rect 80270 -87864 80328 -87854
rect 76832 -89036 76890 -89026
rect 77010 -87890 77014 -87880
rect 77010 -89036 77072 -89026
rect 77188 -87880 77246 -87870
rect 77188 -89042 77246 -89032
rect 77368 -87878 77426 -87868
rect 77368 -89040 77426 -89030
rect 77542 -87878 77600 -87868
rect 77542 -89040 77600 -89030
rect 77720 -87874 77778 -87864
rect 80270 -89026 80328 -89016
rect 80450 -87860 80508 -87850
rect 80450 -89022 80508 -89012
rect 80638 -87860 80696 -87850
rect 80818 -87856 80852 -87850
rect 80996 -87854 81030 -87850
rect 80638 -89022 80696 -89012
rect 80812 -87866 80870 -87856
rect 80462 -89026 80496 -89022
rect 80640 -89026 80674 -89022
rect 77720 -89036 77778 -89026
rect 80812 -89028 80870 -89018
rect 80988 -87864 81046 -87854
rect 81174 -87856 81208 -87850
rect 81352 -87856 81386 -87850
rect 81530 -87854 81564 -87850
rect 81708 -87854 81742 -87850
rect 80988 -89018 80990 -89016
rect 81042 -89018 81046 -89016
rect 80988 -89026 81046 -89018
rect 81170 -87866 81228 -87856
rect 81348 -87866 81406 -87856
rect 80990 -89028 81042 -89026
rect 81170 -89028 81228 -89018
rect 81346 -87882 81348 -87872
rect 81346 -89028 81406 -89018
rect 81522 -87864 81580 -87854
rect 81522 -89026 81580 -89016
rect 81702 -87864 81760 -87854
rect 81886 -87856 81920 -87850
rect 81702 -89026 81760 -89016
rect 81876 -87866 81934 -87856
rect 82064 -87860 82098 -87850
rect 81876 -89028 81934 -89018
rect 82058 -87870 82116 -87860
rect 82242 -87862 82276 -87850
rect 82420 -87854 82454 -87850
rect 82058 -89032 82116 -89022
rect 82232 -87872 82290 -87862
rect 82232 -89034 82290 -89024
rect 82410 -87864 82468 -87854
rect 82598 -87860 82632 -87850
rect 82776 -87860 82810 -87850
rect 82954 -87858 82988 -87850
rect 83132 -87858 83166 -87850
rect 82410 -89026 82468 -89016
rect 82592 -87870 82650 -87860
rect 82592 -89032 82650 -89022
rect 82766 -87870 82824 -87860
rect 82766 -89032 82824 -89022
rect 82946 -87868 83004 -87858
rect 83128 -87868 83186 -87858
rect 83310 -87864 83344 -87850
rect 83488 -87862 83522 -87850
rect 83666 -87862 83700 -87850
rect 83844 -87858 83878 -87850
rect 82946 -89030 83004 -89020
rect 83124 -87884 83128 -87874
rect 83124 -89030 83186 -89020
rect 83302 -87874 83360 -87864
rect 83302 -89036 83360 -89026
rect 83482 -87872 83540 -87862
rect 83482 -89034 83540 -89024
rect 83656 -87872 83714 -87862
rect 83656 -89034 83714 -89024
rect 83834 -87868 83892 -87858
rect 83834 -89030 83892 -89020
rect 68330 -89073 68424 -89072
rect 68510 -89073 68604 -89072
rect 68690 -89073 68784 -89072
rect 68868 -89073 68962 -89072
rect 69044 -89073 69138 -89072
rect 69400 -89073 69494 -89072
rect 69578 -89073 69672 -89072
rect 69760 -89073 69854 -89072
rect 69934 -89073 70028 -89070
rect 70114 -89073 70208 -89072
rect 70470 -89073 70564 -89072
rect 70644 -89073 70738 -89070
rect 70824 -89073 70918 -89068
rect 71002 -89073 71096 -89072
rect 71180 -89073 71274 -89070
rect 71360 -89073 71454 -89072
rect 71536 -89073 71630 -89072
rect 71714 -89073 71808 -89072
rect 74226 -89073 74320 -89070
rect 74406 -89073 74500 -89070
rect 74586 -89073 74680 -89070
rect 74764 -89073 74858 -89070
rect 74940 -89073 75034 -89070
rect 75120 -89073 75214 -89072
rect 75296 -89073 75390 -89070
rect 75474 -89073 75568 -89070
rect 75656 -89073 75750 -89070
rect 75830 -89073 75924 -89068
rect 76010 -89073 76104 -89070
rect 76186 -89073 76280 -89072
rect 76366 -89073 76460 -89070
rect 76540 -89073 76634 -89068
rect 76720 -89073 76814 -89066
rect 76898 -89073 76992 -89070
rect 77076 -89073 77170 -89068
rect 77256 -89073 77350 -89070
rect 77432 -89073 77526 -89070
rect 77610 -89073 77704 -89070
rect 80340 -89073 80434 -89064
rect 80520 -89073 80614 -89064
rect 80700 -89073 80794 -89064
rect 80878 -89073 80972 -89064
rect 81054 -89073 81148 -89064
rect 81234 -89073 81328 -89066
rect 81410 -89073 81504 -89064
rect 81588 -89073 81682 -89064
rect 81770 -89073 81864 -89064
rect 81944 -89072 82038 -89062
rect 68330 -89074 81944 -89073
rect 66107 -89076 80340 -89074
rect 66107 -89078 76720 -89076
rect 66107 -89080 70824 -89078
rect 66107 -89082 69934 -89080
rect 56390 -89192 64384 -89126
rect 56390 -89246 56418 -89192
rect 56534 -89194 56968 -89192
rect 56534 -89246 56598 -89194
rect 56390 -89248 56598 -89246
rect 56714 -89248 56784 -89194
rect 56900 -89246 56968 -89194
rect 57084 -89246 57144 -89192
rect 57260 -89246 57318 -89192
rect 57434 -89194 64384 -89192
rect 57434 -89246 57494 -89194
rect 56900 -89248 57494 -89246
rect 57610 -89196 64384 -89194
rect 57610 -89200 61594 -89196
rect 57610 -89248 57682 -89200
rect 56390 -89254 57682 -89248
rect 57798 -89254 57856 -89200
rect 57972 -89204 61594 -89200
rect 57972 -89208 59468 -89204
rect 57972 -89210 58412 -89208
rect 57972 -89212 58214 -89210
rect 57972 -89254 58038 -89212
rect 56390 -89258 58038 -89254
rect 56362 -89326 56416 -89306
rect 56414 -90484 56416 -89326
rect 56546 -89316 56582 -89258
rect 56546 -89326 56600 -89316
rect 56546 -89328 56548 -89326
rect 56542 -89338 56548 -89328
rect 56708 -89324 56762 -89306
rect 56908 -89316 56944 -89258
rect 57068 -89316 57122 -89306
rect 57260 -89316 57296 -89258
rect 56600 -89338 56602 -89328
rect 56542 -90482 56548 -90472
rect 56362 -91031 56416 -90484
rect 56546 -90484 56548 -90482
rect 56600 -90482 56602 -90472
rect 56708 -89334 56772 -89324
rect 56906 -89326 56958 -89316
rect 57068 -89326 57124 -89316
rect 56546 -90486 56600 -90484
rect 56548 -90494 56600 -90486
rect 56708 -90492 56720 -89334
rect 56900 -89336 56906 -89326
rect 56958 -89336 56960 -89326
rect 56900 -90480 56906 -90470
rect 56708 -90502 56772 -90492
rect 56958 -90480 56960 -90470
rect 56906 -90494 56958 -90484
rect 57068 -90484 57072 -89326
rect 57260 -89326 57312 -89316
rect 57068 -90494 57124 -90484
rect 57254 -89342 57260 -89332
rect 57426 -89318 57480 -89306
rect 57616 -89316 57652 -89258
rect 57682 -89264 57798 -89258
rect 57856 -89264 58006 -89258
rect 57616 -89318 57656 -89316
rect 57426 -89328 57486 -89318
rect 57312 -89342 57314 -89332
rect 57254 -90484 57260 -90476
rect 57312 -90484 57314 -90476
rect 57254 -90486 57314 -90484
rect 57426 -90486 57434 -89328
rect 57614 -89328 57666 -89318
rect 57260 -90494 57312 -90486
rect 56708 -90540 56762 -90502
rect 56710 -91031 56758 -90540
rect 57068 -91031 57122 -90494
rect 57426 -90496 57486 -90486
rect 57608 -89348 57614 -89338
rect 57780 -89328 57834 -89306
rect 57666 -89348 57668 -89338
rect 57608 -90486 57614 -90482
rect 57666 -90486 57668 -90482
rect 57608 -90492 57668 -90486
rect 57832 -90486 57834 -89328
rect 57970 -89316 58006 -89264
rect 58154 -89258 58214 -89212
rect 58038 -89276 58154 -89266
rect 58292 -89258 58412 -89210
rect 58214 -89278 58292 -89268
rect 58136 -89308 58190 -89306
rect 57970 -89326 58026 -89316
rect 57970 -89334 57974 -89326
rect 57614 -90496 57666 -90492
rect 57426 -91031 57480 -90496
rect 57780 -91031 57834 -90486
rect 57964 -89344 57974 -89334
rect 57964 -90484 57974 -90478
rect 57964 -90488 58026 -90484
rect 57974 -90494 58026 -90488
rect 58136 -89318 58194 -89308
rect 58332 -89312 58368 -89258
rect 58490 -89258 58574 -89208
rect 58412 -89276 58490 -89266
rect 58652 -89258 58760 -89208
rect 58574 -89276 58652 -89266
rect 58136 -90476 58142 -89318
rect 58328 -89322 58380 -89312
rect 58136 -90486 58194 -90476
rect 58322 -89340 58328 -89330
rect 58494 -89316 58548 -89306
rect 58684 -89312 58720 -89258
rect 58838 -89210 59108 -89208
rect 58838 -89258 58936 -89210
rect 58760 -89276 58838 -89266
rect 59014 -89258 59108 -89210
rect 58936 -89278 59014 -89268
rect 58494 -89326 58552 -89316
rect 58684 -89322 58738 -89312
rect 58684 -89324 58686 -89322
rect 58380 -89340 58382 -89330
rect 58322 -90480 58328 -90474
rect 58380 -90480 58382 -90474
rect 58322 -90484 58382 -90480
rect 58494 -90484 58500 -89326
rect 58682 -89334 58686 -89324
rect 58852 -89316 58906 -89306
rect 58738 -89334 58742 -89324
rect 58682 -90478 58686 -90468
rect 58136 -91031 58190 -90486
rect 58328 -90490 58380 -90484
rect 58334 -90492 58368 -90490
rect 58494 -90494 58552 -90484
rect 58738 -90478 58742 -90468
rect 58852 -89326 58910 -89316
rect 59044 -89318 59080 -89258
rect 59186 -89258 59292 -89208
rect 59108 -89276 59186 -89266
rect 59370 -89258 59468 -89208
rect 59292 -89276 59370 -89266
rect 58686 -90490 58738 -90480
rect 58852 -90484 58858 -89326
rect 59038 -89328 59090 -89318
rect 58690 -90492 58724 -90490
rect 58852 -90494 58910 -90484
rect 59028 -89346 59038 -89336
rect 59028 -90486 59038 -90480
rect 59028 -90490 59090 -90486
rect 58494 -91031 58548 -90494
rect 58852 -91031 58906 -90494
rect 59038 -90496 59090 -90490
rect 59208 -89320 59262 -89306
rect 59402 -89318 59438 -89258
rect 59546 -89258 59642 -89204
rect 59468 -89272 59546 -89262
rect 59720 -89208 60874 -89204
rect 59720 -89258 59832 -89208
rect 59642 -89272 59720 -89262
rect 59558 -89316 59612 -89306
rect 59750 -89316 59786 -89258
rect 59910 -89258 60874 -89208
rect 59832 -89276 59910 -89266
rect 60952 -89208 61416 -89204
rect 60952 -89258 61064 -89208
rect 60874 -89272 60952 -89262
rect 61142 -89210 61416 -89208
rect 61142 -89258 61242 -89210
rect 61064 -89276 61142 -89266
rect 61320 -89258 61416 -89210
rect 61242 -89278 61320 -89268
rect 61494 -89254 61594 -89204
rect 61672 -89200 64384 -89196
rect 61672 -89204 62122 -89200
rect 61672 -89254 61770 -89204
rect 61494 -89258 61770 -89254
rect 61416 -89272 61494 -89262
rect 61594 -89264 61672 -89258
rect 61848 -89258 61962 -89204
rect 61770 -89272 61848 -89262
rect 62040 -89258 62122 -89204
rect 62200 -89204 62842 -89200
rect 62200 -89258 62298 -89204
rect 61962 -89272 62040 -89262
rect 62122 -89268 62200 -89258
rect 62376 -89258 62478 -89204
rect 62298 -89272 62376 -89262
rect 62556 -89208 62842 -89204
rect 62556 -89258 62652 -89208
rect 62478 -89272 62556 -89262
rect 62730 -89258 62842 -89208
rect 62920 -89258 63026 -89200
rect 63104 -89258 63188 -89200
rect 63266 -89204 63716 -89200
rect 63266 -89258 63370 -89204
rect 62652 -89276 62730 -89266
rect 62842 -89268 62920 -89258
rect 63026 -89268 63104 -89258
rect 63188 -89268 63266 -89258
rect 63448 -89208 63716 -89204
rect 63448 -89258 63554 -89208
rect 63370 -89272 63448 -89262
rect 63632 -89258 63716 -89208
rect 63794 -89258 63900 -89200
rect 63978 -89258 64088 -89200
rect 64166 -89258 64256 -89200
rect 64334 -89258 64384 -89200
rect 66107 -89227 68330 -89082
rect 63554 -89276 63632 -89266
rect 63716 -89268 63794 -89258
rect 63900 -89268 63978 -89258
rect 64088 -89268 64166 -89258
rect 64256 -89268 64334 -89258
rect 60802 -89306 60838 -89304
rect 61166 -89306 61202 -89304
rect 62584 -89306 62620 -89302
rect 63304 -89306 63340 -89304
rect 63652 -89306 63688 -89304
rect 64008 -89306 64044 -89302
rect 59916 -89312 59970 -89306
rect 59208 -89330 59266 -89320
rect 59396 -89328 59448 -89318
rect 59208 -90488 59214 -89330
rect 59388 -89338 59396 -89328
rect 59388 -90482 59396 -90472
rect 59208 -90498 59266 -90488
rect 59396 -90496 59448 -90486
rect 59558 -89326 59622 -89316
rect 59750 -89320 59804 -89316
rect 59558 -90484 59570 -89326
rect 59746 -89326 59806 -89320
rect 59746 -89330 59752 -89326
rect 59804 -89330 59806 -89326
rect 59746 -90474 59752 -90464
rect 59750 -90478 59752 -90474
rect 59558 -90494 59622 -90484
rect 59804 -90474 59806 -90464
rect 59916 -89322 59974 -89312
rect 59752 -90494 59804 -90484
rect 59916 -90480 59922 -89322
rect 59916 -90490 59974 -90480
rect 60794 -89326 60848 -89306
rect 60794 -90484 60796 -89326
rect 60980 -89326 61032 -89316
rect 60974 -89340 60980 -89330
rect 61140 -89326 61202 -89306
rect 61500 -89310 61554 -89306
rect 61340 -89318 61374 -89316
rect 61032 -89340 61034 -89330
rect 60974 -90484 60980 -90474
rect 61032 -90484 61034 -90474
rect 61140 -90484 61142 -89326
rect 61194 -90484 61202 -89326
rect 61330 -89328 61382 -89318
rect 59208 -90540 59262 -90498
rect 59210 -91031 59262 -90540
rect 59558 -91031 59612 -90494
rect 59916 -91031 59970 -90490
rect 60794 -90495 60848 -90484
rect 60980 -90494 61032 -90484
rect 60802 -91031 60838 -90495
rect 61140 -91031 61202 -90484
rect 61322 -89342 61330 -89332
rect 61322 -90486 61330 -90476
rect 61330 -90496 61382 -90486
rect 61500 -89328 61560 -89310
rect 61696 -89318 61730 -89316
rect 61690 -89324 61742 -89318
rect 61500 -90486 61506 -89328
rect 61558 -90486 61560 -89328
rect 61680 -89328 61742 -89324
rect 61680 -89334 61690 -89328
rect 61680 -90478 61690 -90468
rect 61500 -91031 61560 -90486
rect 61690 -90496 61742 -90486
rect 61858 -89322 61912 -89306
rect 62212 -89312 62266 -89306
rect 61858 -89332 61914 -89322
rect 61858 -90490 61862 -89332
rect 61858 -90495 61914 -90490
rect 62042 -89326 62094 -89316
rect 62212 -89322 62268 -89312
rect 62094 -89344 62102 -89334
rect 62094 -90484 62102 -90478
rect 62042 -90488 62102 -90484
rect 62212 -90480 62216 -89322
rect 62268 -90480 62272 -89324
rect 62398 -89326 62450 -89316
rect 62042 -90494 62094 -90488
rect 62212 -90495 62272 -90480
rect 62396 -89348 62398 -89338
rect 62568 -89322 62622 -89306
rect 62926 -89312 62980 -89306
rect 62450 -89348 62456 -89338
rect 62396 -90484 62398 -90482
rect 62450 -90484 62456 -90482
rect 62396 -90492 62456 -90484
rect 62568 -90480 62570 -89322
rect 62756 -89326 62808 -89316
rect 62398 -90494 62450 -90492
rect 61862 -90500 61914 -90495
rect 61862 -91031 61912 -90500
rect 62220 -91031 62272 -90495
rect 62568 -90497 62622 -90480
rect 62752 -89348 62756 -89338
rect 62926 -89326 62984 -89312
rect 62808 -89348 62812 -89338
rect 62752 -90484 62756 -90482
rect 62808 -90484 62812 -90482
rect 62752 -90492 62812 -90484
rect 62978 -90484 62984 -89326
rect 63112 -89320 63164 -89310
rect 63106 -89340 63112 -89330
rect 63284 -89322 63340 -89306
rect 63476 -89318 63510 -89316
rect 63164 -89340 63166 -89330
rect 63106 -90478 63112 -90474
rect 63164 -90478 63166 -90474
rect 63106 -90484 63166 -90478
rect 63284 -90480 63288 -89322
rect 63468 -89328 63520 -89318
rect 63640 -89322 63694 -89306
rect 62756 -90494 62808 -90492
rect 62573 -91031 62620 -90497
rect 62926 -91031 62984 -90484
rect 63112 -90488 63164 -90484
rect 63120 -90492 63154 -90488
rect 63284 -91031 63340 -90480
rect 63466 -89352 63468 -89342
rect 63638 -89332 63694 -89322
rect 63520 -89352 63526 -89342
rect 63466 -90496 63526 -90486
rect 63690 -90490 63694 -89332
rect 63638 -90497 63694 -90490
rect 63826 -89326 63878 -89316
rect 63990 -89318 64044 -89306
rect 63990 -89328 64046 -89318
rect 63878 -89344 63886 -89334
rect 63878 -90484 63886 -90478
rect 63826 -90488 63886 -90484
rect 63990 -90486 63994 -89328
rect 64184 -89326 64236 -89316
rect 63826 -90494 63878 -90488
rect 63990 -90496 64046 -90486
rect 64182 -89348 64184 -89338
rect 64348 -89328 64402 -89306
rect 64236 -89348 64242 -89338
rect 64182 -90484 64184 -90482
rect 64236 -90484 64242 -90482
rect 64182 -90492 64242 -90484
rect 64400 -90486 64402 -89328
rect 64184 -90494 64236 -90492
rect 63638 -90500 63690 -90497
rect 63638 -91031 63688 -90500
rect 63990 -91031 64044 -90496
rect 64348 -91031 64402 -90486
rect 65342 -89783 65498 -89782
rect 67554 -89783 67842 -89227
rect 68424 -89227 68510 -89082
rect 68330 -89238 68424 -89228
rect 68604 -89227 68690 -89082
rect 68510 -89238 68604 -89228
rect 68784 -89227 68868 -89082
rect 68690 -89238 68784 -89228
rect 68962 -89227 69044 -89082
rect 68868 -89238 68962 -89228
rect 69138 -89084 69400 -89082
rect 69138 -89227 69224 -89084
rect 69044 -89238 69138 -89228
rect 69318 -89227 69400 -89084
rect 69224 -89240 69318 -89230
rect 69494 -89227 69578 -89082
rect 69400 -89238 69494 -89228
rect 69672 -89227 69760 -89082
rect 69578 -89238 69672 -89228
rect 69854 -89226 69934 -89082
rect 70028 -89082 70644 -89080
rect 70028 -89226 70114 -89082
rect 69854 -89227 70114 -89226
rect 69760 -89238 69854 -89228
rect 69934 -89236 70028 -89227
rect 70208 -89084 70470 -89082
rect 70208 -89227 70290 -89084
rect 70114 -89238 70208 -89228
rect 70384 -89227 70470 -89084
rect 70290 -89240 70384 -89230
rect 70564 -89226 70644 -89082
rect 70738 -89224 70824 -89080
rect 70918 -89080 75830 -89078
rect 70918 -89082 71180 -89080
rect 70918 -89224 71002 -89082
rect 70738 -89226 71002 -89224
rect 70564 -89227 71002 -89226
rect 70470 -89238 70564 -89228
rect 70644 -89236 70738 -89227
rect 70824 -89234 70918 -89227
rect 71096 -89226 71180 -89082
rect 71274 -89082 74226 -89080
rect 71274 -89226 71360 -89082
rect 71096 -89227 71360 -89226
rect 71002 -89238 71096 -89228
rect 71180 -89236 71274 -89227
rect 71454 -89227 71536 -89082
rect 71360 -89238 71454 -89228
rect 71630 -89227 71714 -89082
rect 71536 -89238 71630 -89228
rect 71808 -89226 74226 -89082
rect 74320 -89226 74406 -89080
rect 74500 -89226 74586 -89080
rect 74680 -89226 74764 -89080
rect 74858 -89226 74940 -89080
rect 75034 -89082 75296 -89080
rect 75034 -89226 75120 -89082
rect 71808 -89227 75120 -89226
rect 71714 -89238 71808 -89228
rect 74226 -89236 74320 -89227
rect 74406 -89236 74500 -89227
rect 74586 -89236 74680 -89227
rect 74764 -89236 74858 -89227
rect 74940 -89236 75034 -89227
rect 75214 -89226 75296 -89082
rect 75390 -89226 75474 -89080
rect 75568 -89226 75656 -89080
rect 75750 -89224 75830 -89080
rect 75924 -89080 76540 -89078
rect 75924 -89224 76010 -89080
rect 75750 -89226 76010 -89224
rect 76104 -89082 76366 -89080
rect 76104 -89226 76186 -89082
rect 75214 -89227 76186 -89226
rect 75120 -89238 75214 -89228
rect 75296 -89236 75390 -89227
rect 75474 -89236 75568 -89227
rect 75656 -89236 75750 -89227
rect 75830 -89234 75924 -89227
rect 76010 -89236 76104 -89227
rect 76280 -89226 76366 -89082
rect 76460 -89224 76540 -89080
rect 76634 -89222 76720 -89078
rect 76814 -89078 80340 -89076
rect 76814 -89080 77076 -89078
rect 76814 -89222 76898 -89080
rect 76634 -89224 76898 -89222
rect 76460 -89226 76898 -89224
rect 76992 -89224 77076 -89080
rect 77170 -89080 80340 -89078
rect 77170 -89224 77256 -89080
rect 76992 -89226 77256 -89224
rect 77350 -89226 77432 -89080
rect 77526 -89226 77610 -89080
rect 77704 -89220 80340 -89080
rect 80434 -89220 80520 -89074
rect 80614 -89220 80700 -89074
rect 80794 -89220 80878 -89074
rect 80972 -89220 81054 -89074
rect 81148 -89076 81410 -89074
rect 81148 -89220 81234 -89076
rect 77704 -89222 81234 -89220
rect 81328 -89220 81410 -89076
rect 81504 -89220 81588 -89074
rect 81682 -89220 81770 -89074
rect 81864 -89218 81944 -89074
rect 82124 -89073 82218 -89064
rect 82300 -89073 82394 -89066
rect 82480 -89073 82574 -89064
rect 82654 -89072 82748 -89062
rect 82038 -89074 82654 -89073
rect 82038 -89218 82124 -89074
rect 81864 -89220 82124 -89218
rect 82218 -89076 82480 -89074
rect 82218 -89220 82300 -89076
rect 81328 -89222 82300 -89220
rect 82394 -89220 82480 -89076
rect 82574 -89218 82654 -89074
rect 82834 -89070 82928 -89060
rect 82748 -89216 82834 -89073
rect 83012 -89073 83106 -89064
rect 83190 -89072 83284 -89062
rect 82928 -89074 83190 -89073
rect 82928 -89216 83012 -89074
rect 82748 -89218 83012 -89216
rect 82574 -89220 83012 -89218
rect 83106 -89218 83190 -89074
rect 83370 -89073 83464 -89064
rect 83546 -89073 83640 -89064
rect 83724 -89073 83818 -89064
rect 83284 -89074 83919 -89073
rect 83284 -89218 83370 -89074
rect 83106 -89220 83370 -89218
rect 83464 -89220 83546 -89074
rect 83640 -89220 83724 -89074
rect 83818 -89220 83919 -89074
rect 82394 -89222 83919 -89220
rect 77704 -89226 83919 -89222
rect 76280 -89227 83919 -89226
rect 76186 -89238 76280 -89228
rect 76366 -89236 76460 -89227
rect 76540 -89234 76634 -89227
rect 76720 -89232 76814 -89227
rect 76898 -89236 76992 -89227
rect 77076 -89234 77170 -89227
rect 77256 -89236 77350 -89227
rect 77432 -89236 77526 -89227
rect 77610 -89236 77704 -89227
rect 80340 -89230 80434 -89227
rect 80520 -89230 80614 -89227
rect 80700 -89230 80794 -89227
rect 80878 -89230 80972 -89227
rect 81054 -89230 81148 -89227
rect 81234 -89232 81328 -89227
rect 81410 -89230 81504 -89227
rect 81588 -89230 81682 -89227
rect 81770 -89230 81864 -89227
rect 81944 -89228 82038 -89227
rect 82124 -89230 82218 -89227
rect 82300 -89232 82394 -89227
rect 82480 -89230 82574 -89227
rect 82654 -89228 82748 -89227
rect 83012 -89230 83106 -89227
rect 83190 -89228 83284 -89227
rect 83370 -89230 83464 -89227
rect 83546 -89230 83640 -89227
rect 83724 -89230 83818 -89227
rect 68274 -89290 68308 -89276
rect 68452 -89284 68486 -89276
rect 68630 -89280 68664 -89276
rect 65342 -90049 67842 -89783
rect 68268 -89300 68326 -89290
rect 65342 -90547 67819 -90049
rect 68268 -90462 68326 -90452
rect 68444 -89294 68502 -89284
rect 68622 -89290 68680 -89280
rect 68808 -89286 68842 -89276
rect 68444 -90456 68502 -90446
rect 68620 -89306 68622 -89296
rect 68620 -90452 68680 -90442
rect 68800 -89296 68858 -89286
rect 68986 -89288 69020 -89276
rect 69164 -89284 69198 -89276
rect 68800 -90458 68858 -90448
rect 68980 -89298 69038 -89288
rect 68980 -90460 69038 -90450
rect 69156 -89294 69214 -89284
rect 69342 -89288 69376 -89276
rect 69520 -89282 69554 -89276
rect 69156 -90456 69214 -90446
rect 69332 -89298 69390 -89288
rect 69332 -90460 69390 -90450
rect 69508 -89292 69566 -89282
rect 69698 -89284 69732 -89276
rect 69508 -90454 69566 -90444
rect 69688 -89294 69746 -89284
rect 69876 -89288 69910 -89276
rect 70054 -89284 70088 -89276
rect 70232 -89282 70266 -89276
rect 69688 -90456 69746 -90446
rect 69864 -89298 69922 -89288
rect 69864 -90460 69922 -90450
rect 70044 -89294 70102 -89284
rect 70044 -90456 70102 -90446
rect 70226 -89292 70284 -89282
rect 70410 -89284 70444 -89276
rect 70588 -89284 70622 -89276
rect 70766 -89284 70800 -89276
rect 70944 -89284 70978 -89276
rect 71122 -89278 71156 -89276
rect 70226 -90454 70284 -90444
rect 70406 -89294 70464 -89284
rect 70406 -90456 70464 -90446
rect 70578 -89294 70636 -89284
rect 70578 -90456 70636 -90446
rect 70756 -89294 70814 -89284
rect 70756 -90456 70814 -90446
rect 70934 -89294 70992 -89284
rect 70934 -90456 70992 -90446
rect 71112 -89288 71170 -89278
rect 71300 -89288 71334 -89276
rect 71294 -89298 71352 -89288
rect 71478 -89290 71512 -89276
rect 71656 -89284 71690 -89276
rect 71112 -90442 71114 -90440
rect 71166 -90442 71170 -90440
rect 71112 -90450 71170 -90442
rect 71292 -89312 71294 -89302
rect 71292 -90450 71294 -90448
rect 71114 -90452 71166 -90450
rect 71292 -90458 71352 -90450
rect 71294 -90460 71352 -90458
rect 71472 -89300 71530 -89290
rect 71472 -90462 71530 -90452
rect 71646 -89294 71704 -89284
rect 71834 -89288 71868 -89276
rect 74170 -89288 74204 -89274
rect 74348 -89282 74382 -89274
rect 74526 -89278 74560 -89274
rect 71646 -90456 71704 -90446
rect 71826 -89298 71884 -89288
rect 71826 -90460 71884 -90450
rect 74164 -89298 74222 -89288
rect 74164 -90460 74222 -90450
rect 74340 -89292 74398 -89282
rect 74518 -89288 74576 -89278
rect 74704 -89284 74738 -89274
rect 74340 -90454 74398 -90444
rect 74516 -89304 74518 -89294
rect 74516 -90450 74576 -90440
rect 74696 -89294 74754 -89284
rect 74882 -89286 74916 -89274
rect 75060 -89282 75094 -89274
rect 74696 -90456 74754 -90446
rect 74876 -89296 74934 -89286
rect 74876 -90458 74934 -90448
rect 75052 -89292 75110 -89282
rect 75238 -89286 75272 -89274
rect 75416 -89280 75450 -89274
rect 75052 -90454 75110 -90444
rect 75228 -89296 75286 -89286
rect 75228 -90458 75286 -90448
rect 75404 -89290 75462 -89280
rect 75594 -89282 75628 -89274
rect 75404 -90452 75462 -90442
rect 75584 -89292 75642 -89282
rect 75772 -89286 75806 -89274
rect 75950 -89282 75984 -89274
rect 76128 -89280 76162 -89274
rect 75584 -90454 75642 -90444
rect 75760 -89296 75818 -89286
rect 75760 -90458 75818 -90448
rect 75940 -89292 75998 -89282
rect 75940 -90454 75998 -90444
rect 76122 -89290 76180 -89280
rect 76306 -89282 76340 -89274
rect 76484 -89282 76518 -89274
rect 76662 -89282 76696 -89274
rect 76840 -89282 76874 -89274
rect 77018 -89276 77052 -89274
rect 76122 -90452 76180 -90442
rect 76302 -89292 76360 -89282
rect 76302 -90454 76360 -90444
rect 76474 -89292 76532 -89282
rect 76474 -90454 76532 -90444
rect 76652 -89292 76710 -89282
rect 76652 -90454 76710 -90444
rect 76830 -89292 76888 -89282
rect 76830 -90454 76888 -90444
rect 77008 -89286 77066 -89276
rect 77196 -89286 77230 -89274
rect 77190 -89296 77248 -89286
rect 77374 -89288 77408 -89274
rect 77552 -89282 77586 -89274
rect 77008 -90440 77010 -90438
rect 77062 -90440 77066 -90438
rect 77008 -90448 77066 -90440
rect 77188 -89310 77190 -89300
rect 77188 -90448 77190 -90446
rect 77010 -90450 77062 -90448
rect 77188 -90456 77248 -90448
rect 77190 -90458 77248 -90456
rect 77368 -89298 77426 -89288
rect 77368 -90460 77426 -90450
rect 77542 -89292 77600 -89282
rect 77730 -89286 77764 -89274
rect 80284 -89282 80318 -89268
rect 80462 -89276 80496 -89268
rect 80640 -89272 80674 -89268
rect 77542 -90454 77600 -90444
rect 77722 -89296 77780 -89286
rect 77722 -90458 77780 -90448
rect 80278 -89292 80336 -89282
rect 80278 -90454 80336 -90444
rect 80454 -89286 80512 -89276
rect 80632 -89282 80690 -89272
rect 80818 -89278 80852 -89268
rect 80454 -90448 80512 -90438
rect 80630 -89298 80632 -89288
rect 80630 -90444 80690 -90434
rect 80810 -89288 80868 -89278
rect 80996 -89280 81030 -89268
rect 81174 -89276 81208 -89268
rect 80810 -90450 80868 -90440
rect 80990 -89290 81048 -89280
rect 80990 -90452 81048 -90442
rect 81166 -89286 81224 -89276
rect 81352 -89280 81386 -89268
rect 81530 -89274 81564 -89268
rect 81166 -90448 81224 -90438
rect 81342 -89290 81400 -89280
rect 81342 -90452 81400 -90442
rect 81518 -89284 81576 -89274
rect 81708 -89276 81742 -89268
rect 81518 -90446 81576 -90436
rect 81698 -89286 81756 -89276
rect 81886 -89280 81920 -89268
rect 82064 -89276 82098 -89268
rect 82242 -89274 82276 -89268
rect 81698 -90448 81756 -90438
rect 81874 -89290 81932 -89280
rect 81874 -90452 81932 -90442
rect 82054 -89286 82112 -89276
rect 82054 -90448 82112 -90438
rect 82236 -89284 82294 -89274
rect 82420 -89276 82454 -89268
rect 82598 -89276 82632 -89268
rect 82776 -89276 82810 -89268
rect 82954 -89276 82988 -89268
rect 83132 -89270 83166 -89268
rect 82236 -90446 82294 -90436
rect 82416 -89286 82474 -89276
rect 82416 -90448 82474 -90438
rect 82588 -89286 82646 -89276
rect 82588 -90448 82646 -90438
rect 82766 -89286 82824 -89276
rect 82766 -90448 82824 -90438
rect 82944 -89286 83002 -89276
rect 82944 -90448 83002 -90438
rect 83122 -89280 83180 -89270
rect 83310 -89280 83344 -89268
rect 83304 -89290 83362 -89280
rect 83488 -89282 83522 -89268
rect 83666 -89276 83700 -89268
rect 83122 -90434 83124 -90432
rect 83176 -90434 83180 -90432
rect 83122 -90442 83180 -90434
rect 83302 -89304 83304 -89294
rect 83302 -90442 83304 -90440
rect 83124 -90444 83176 -90442
rect 83302 -90450 83362 -90442
rect 83304 -90452 83362 -90450
rect 83482 -89292 83540 -89282
rect 83482 -90454 83540 -90444
rect 83656 -89286 83714 -89276
rect 83844 -89280 83878 -89268
rect 83656 -90448 83714 -90438
rect 83836 -89290 83894 -89280
rect 83836 -90452 83894 -90442
rect 54869 -91122 86347 -91031
rect 54869 -91190 86365 -91122
rect 54869 -91892 55054 -91190
rect 85992 -91511 86365 -91190
rect 85992 -91728 86360 -91511
rect 85992 -91892 86347 -91728
rect 54869 -91946 86347 -91892
<< via2 >>
rect 60946 -71284 60954 -70134
rect 60954 -71284 61012 -70134
rect 61012 -71284 61016 -70134
rect 61302 -71286 61310 -70138
rect 61310 -71286 61368 -70138
rect 61368 -71286 61372 -70138
rect 61302 -71288 61372 -71286
rect 61654 -71286 61664 -70142
rect 61664 -71286 61722 -70142
rect 61722 -71286 61724 -70142
rect 61654 -71292 61724 -71286
rect 62004 -71280 62022 -70130
rect 62022 -71280 62074 -70130
rect 62366 -71286 62376 -70144
rect 62376 -71286 62434 -70144
rect 62434 -71286 62436 -70144
rect 62366 -71294 62436 -71286
rect 62726 -71284 62730 -70142
rect 62730 -71284 62788 -70142
rect 62788 -71284 62796 -70142
rect 62726 -71292 62796 -71284
rect 63088 -71280 63090 -70130
rect 63090 -71280 63148 -70130
rect 63148 -71280 63158 -70130
rect 63436 -70132 63506 -70130
rect 63436 -71280 63446 -70132
rect 63446 -71280 63504 -70132
rect 63504 -71280 63506 -70132
rect 63794 -70130 63864 -70128
rect 63794 -71278 63802 -70130
rect 63802 -71278 63860 -70130
rect 63860 -71278 63864 -70130
rect 64150 -70130 64220 -70124
rect 64150 -71274 64160 -70130
rect 64160 -71274 64218 -70130
rect 64218 -71274 64220 -70130
rect 68320 -70128 68382 -70126
rect 68320 -71270 68374 -70128
rect 68374 -71270 68382 -70128
rect 68670 -70124 68732 -70122
rect 68670 -71266 68724 -70124
rect 68724 -71266 68732 -70124
rect 69026 -70118 69088 -70116
rect 69026 -71260 69080 -70118
rect 69080 -71260 69088 -70118
rect 69378 -70122 69440 -70120
rect 69378 -71264 69432 -70122
rect 69432 -71264 69440 -70122
rect 69732 -70120 69794 -70118
rect 69732 -71262 69786 -70120
rect 69786 -71262 69794 -70120
rect 70094 -70124 70156 -70122
rect 70094 -71266 70148 -70124
rect 70148 -71266 70156 -70124
rect 70452 -70116 70514 -70114
rect 70452 -71258 70506 -70116
rect 70506 -71258 70514 -70116
rect 70804 -70112 70866 -70110
rect 70804 -71254 70858 -70112
rect 70858 -71254 70866 -70112
rect 71158 -70116 71220 -70114
rect 71158 -71258 71212 -70116
rect 71212 -71258 71220 -70116
rect 71512 -70116 71574 -70114
rect 71512 -71258 71566 -70116
rect 71566 -71258 71574 -70116
rect 71874 -70116 71936 -70114
rect 71874 -71258 71928 -70116
rect 71928 -71258 71936 -70116
rect 72228 -70120 72290 -70118
rect 72228 -71262 72282 -70120
rect 72282 -71262 72290 -70120
rect 72586 -70120 72648 -70118
rect 72586 -71262 72640 -70120
rect 72640 -71262 72648 -70120
rect 72942 -70116 73004 -70114
rect 72942 -71258 72996 -70116
rect 72996 -71258 73004 -70116
rect 73302 -70116 73364 -70114
rect 73302 -71258 73356 -70116
rect 73356 -71258 73364 -70116
rect 73652 -70120 73714 -70118
rect 73652 -71262 73706 -70120
rect 73706 -71262 73714 -70120
rect 74008 -70116 74070 -70114
rect 74008 -71258 74062 -70116
rect 74062 -71258 74070 -70116
rect 74366 -70114 74428 -70112
rect 74366 -71256 74420 -70114
rect 74420 -71256 74428 -70114
rect 74724 -70116 74786 -70114
rect 74724 -71258 74778 -70116
rect 74778 -71258 74786 -70116
rect 75074 -70116 75136 -70114
rect 75074 -71258 75128 -70116
rect 75128 -71258 75136 -70116
rect 75432 -70114 75494 -70112
rect 75432 -71256 75486 -70114
rect 75486 -71256 75494 -70114
rect 75788 -70114 75850 -70112
rect 75788 -71256 75842 -70114
rect 75842 -71256 75850 -70114
rect 76146 -70116 76208 -70114
rect 76146 -71258 76200 -70116
rect 76200 -71258 76208 -70116
rect 76496 -70114 76558 -70112
rect 76496 -71256 76550 -70114
rect 76550 -71256 76558 -70114
rect 76860 -70116 76922 -70114
rect 76860 -71258 76914 -70116
rect 76914 -71258 76922 -70116
rect 77212 -70120 77274 -70118
rect 77212 -71262 77266 -70120
rect 77266 -71262 77274 -70120
rect 77568 -70114 77630 -70112
rect 77568 -71256 77622 -70114
rect 77622 -71256 77630 -70114
rect 77926 -70112 77988 -70110
rect 77926 -71254 77980 -70112
rect 77980 -71254 77988 -70112
rect 78282 -70114 78344 -70112
rect 78282 -71256 78336 -70114
rect 78336 -71256 78344 -70114
rect 78638 -70114 78700 -70112
rect 78638 -71256 78692 -70114
rect 78692 -71256 78700 -70114
rect 78996 -70116 79058 -70114
rect 78996 -71258 79050 -70116
rect 79050 -71258 79058 -70116
rect 79346 -70120 79408 -70118
rect 79346 -71262 79400 -70120
rect 79400 -71262 79408 -70120
rect 79704 -70120 79766 -70118
rect 79704 -71262 79758 -70120
rect 79758 -71262 79766 -70120
rect 80058 -70114 80120 -70112
rect 80058 -71256 80112 -70114
rect 80112 -71256 80120 -70114
rect 80412 -70120 80474 -70118
rect 80412 -71262 80466 -70120
rect 80466 -71262 80474 -70120
rect 80768 -70116 80830 -70114
rect 80768 -71258 80822 -70116
rect 80822 -71258 80830 -70116
rect 81126 -70120 81188 -70118
rect 81126 -71262 81180 -70120
rect 81180 -71262 81188 -70120
rect 81480 -70116 81542 -70114
rect 81480 -71258 81534 -70116
rect 81534 -71258 81542 -70116
rect 81836 -70120 81898 -70118
rect 81836 -71262 81890 -70120
rect 81890 -71262 81898 -70120
rect 82190 -70116 82252 -70114
rect 82190 -71258 82244 -70116
rect 82244 -71258 82252 -70116
rect 82546 -70120 82608 -70118
rect 82546 -71262 82600 -70120
rect 82600 -71262 82608 -70120
rect 82906 -70116 82968 -70114
rect 82906 -71258 82960 -70116
rect 82960 -71258 82968 -70116
rect 83264 -70114 83326 -70112
rect 83264 -71256 83318 -70114
rect 83318 -71256 83326 -70114
rect 83620 -70120 83682 -70118
rect 83620 -71262 83674 -70120
rect 83674 -71262 83682 -70120
rect 83976 -70120 84038 -70118
rect 83976 -71262 84030 -70120
rect 84030 -71262 84038 -70120
rect 68314 -72706 68372 -71562
rect 68372 -72706 68376 -71562
rect 68664 -71554 68726 -71540
rect 68664 -72684 68668 -71554
rect 68668 -72684 68726 -71554
rect 69018 -71554 69080 -71542
rect 69018 -72652 69028 -71554
rect 69028 -72652 69080 -71554
rect 69378 -71558 69440 -71540
rect 69378 -72684 69382 -71558
rect 69382 -72684 69440 -71558
rect 69724 -71562 69786 -71548
rect 69724 -72658 69740 -71562
rect 69740 -72658 69786 -71562
rect 70086 -71560 70148 -71536
rect 70086 -72646 70092 -71560
rect 70092 -72646 70148 -71560
rect 70450 -71560 70512 -71542
rect 70450 -72652 70502 -71560
rect 70502 -72652 70512 -71560
rect 70790 -71560 70852 -71546
rect 70790 -72656 70800 -71560
rect 70800 -72656 70852 -71560
rect 71148 -71558 71210 -71554
rect 71148 -72664 71156 -71558
rect 71156 -72664 71210 -71558
rect 71504 -71558 71566 -71546
rect 71504 -72656 71516 -71558
rect 71516 -72656 71566 -71558
rect 71858 -71558 71920 -71542
rect 71858 -72652 71870 -71558
rect 71870 -72652 71920 -71558
rect 72216 -71558 72278 -71546
rect 72216 -72656 72230 -71558
rect 72230 -72656 72278 -71558
rect 72570 -71560 72632 -71544
rect 72570 -72654 72586 -71560
rect 72586 -72654 72632 -71560
rect 72946 -71558 73008 -71542
rect 72946 -72652 72996 -71558
rect 72996 -72652 73008 -71558
rect 73286 -71562 73348 -71558
rect 73286 -72668 73292 -71562
rect 73292 -72668 73348 -71562
rect 73642 -71560 73704 -71550
rect 73642 -72660 73654 -71560
rect 73654 -72660 73704 -71560
rect 73988 -71554 74050 -71542
rect 73988 -72652 74010 -71554
rect 74010 -72652 74050 -71554
rect 74352 -72670 74364 -71560
rect 74364 -72670 74414 -71560
rect 74714 -72666 74720 -71556
rect 74720 -72666 74776 -71556
rect 75068 -72682 75078 -71572
rect 75078 -72682 75130 -71572
rect 75426 -72670 75432 -71560
rect 75432 -72670 75488 -71560
rect 75764 -71564 75826 -71544
rect 75764 -72654 75786 -71564
rect 75786 -72654 75826 -71564
rect 76130 -71556 76192 -71542
rect 76130 -72652 76146 -71556
rect 76146 -72652 76192 -71556
rect 76478 -71556 76540 -71542
rect 76478 -72652 76500 -71556
rect 76500 -72652 76540 -71556
rect 76854 -71562 76916 -71546
rect 76854 -72656 76912 -71562
rect 76912 -72656 76916 -71562
rect 77196 -71562 77258 -71550
rect 77196 -72660 77212 -71562
rect 77212 -72660 77258 -71562
rect 77548 -72672 77566 -71562
rect 77566 -72672 77610 -71562
rect 77908 -71564 77970 -71538
rect 77908 -72648 77924 -71564
rect 77924 -72648 77970 -71564
rect 78274 -71568 78336 -71540
rect 78274 -72650 78276 -71568
rect 78276 -72650 78334 -71568
rect 78334 -72650 78336 -71568
rect 78624 -71568 78686 -71562
rect 78624 -72672 78636 -71568
rect 78636 -72672 78686 -71568
rect 78990 -71568 79052 -71562
rect 78990 -72672 79048 -71568
rect 79048 -72672 79052 -71568
rect 79338 -71566 79400 -71542
rect 79338 -72652 79344 -71566
rect 79344 -72652 79400 -71566
rect 79692 -71562 79754 -71550
rect 79692 -72660 79700 -71562
rect 79700 -72660 79754 -71562
rect 80048 -71560 80110 -71556
rect 80048 -72666 80058 -71560
rect 80058 -72666 80110 -71560
rect 80398 -72670 80416 -71560
rect 80416 -72670 80460 -71560
rect 80760 -71562 80822 -71552
rect 80760 -72662 80772 -71562
rect 80772 -72662 80822 -71562
rect 81120 -72672 81124 -71562
rect 81124 -72672 81182 -71562
rect 81478 -71556 81540 -71550
rect 81478 -72660 81482 -71556
rect 81482 -72660 81540 -71556
rect 81848 -71556 81910 -71552
rect 81848 -72662 81894 -71556
rect 81894 -72662 81910 -71556
rect 82186 -72670 82196 -71560
rect 82196 -72670 82248 -71560
rect 82542 -72676 82556 -71566
rect 82556 -72676 82604 -71566
rect 82910 -72684 82966 -71574
rect 82966 -72684 82972 -71574
rect 83258 -71554 83320 -71552
rect 83258 -72662 83262 -71554
rect 83262 -72662 83320 -71554
rect 83612 -72684 83622 -71574
rect 83622 -72684 83674 -71574
rect 83962 -71556 84024 -71550
rect 83962 -72660 83978 -71556
rect 83978 -72660 84024 -71556
rect 56488 -74540 56490 -73402
rect 56490 -74540 56544 -73402
rect 56852 -74534 56906 -73396
rect 56906 -74534 56908 -73396
rect 57196 -74546 57202 -73408
rect 57202 -74546 57252 -73408
rect 57556 -74540 57558 -73402
rect 57558 -74540 57612 -73402
rect 57916 -74546 57970 -73408
rect 57970 -74546 57972 -73408
rect 58274 -74548 58276 -73410
rect 58276 -74548 58330 -73410
rect 58628 -73402 58684 -73400
rect 58628 -74538 58630 -73402
rect 58630 -74538 58684 -73402
rect 58980 -74542 58986 -73404
rect 58986 -74542 59036 -73404
rect 59342 -74538 59344 -73400
rect 59344 -74538 59398 -73400
rect 59694 -74542 59698 -73404
rect 59698 -74542 59750 -73404
rect 60052 -74550 60054 -73412
rect 60054 -74550 60108 -73412
rect 60402 -74548 60406 -73410
rect 60406 -74548 60458 -73410
rect 60764 -74544 60768 -73406
rect 60768 -74544 60820 -73406
rect 61118 -74548 61122 -73410
rect 61122 -74548 61174 -73410
rect 61476 -74542 61478 -73404
rect 61478 -74542 61532 -73404
rect 61826 -74548 61828 -73410
rect 61828 -74548 61882 -73410
rect 62188 -74550 62242 -73414
rect 62242 -74550 62244 -73414
rect 62188 -74552 62244 -74550
rect 62544 -74548 62546 -73410
rect 62546 -74548 62600 -73410
rect 62894 -74550 62898 -73414
rect 62898 -74550 62950 -73414
rect 62894 -74552 62950 -74550
rect 63254 -74544 63256 -73412
rect 63256 -74544 63310 -73412
rect 63254 -74550 63310 -74544
rect 63614 -74546 63666 -73414
rect 63666 -74546 63670 -73414
rect 63614 -74552 63670 -74546
rect 63966 -74544 63968 -73408
rect 63968 -74544 64022 -73408
rect 63966 -74546 64022 -74544
rect 64320 -74546 64322 -73408
rect 64322 -74546 64376 -73408
rect 56472 -76002 56474 -74864
rect 56474 -76002 56528 -74864
rect 56836 -75996 56890 -74858
rect 56890 -75996 56892 -74858
rect 57180 -76008 57186 -74870
rect 57186 -76008 57236 -74870
rect 57540 -76002 57542 -74864
rect 57542 -76002 57596 -74864
rect 57900 -76008 57954 -74870
rect 57954 -76008 57956 -74870
rect 58258 -76010 58260 -74872
rect 58260 -76010 58314 -74872
rect 58612 -74864 58668 -74862
rect 58612 -76000 58614 -74864
rect 58614 -76000 58668 -74864
rect 58964 -76004 58970 -74866
rect 58970 -76004 59020 -74866
rect 59326 -76000 59328 -74862
rect 59328 -76000 59382 -74862
rect 59678 -76004 59682 -74866
rect 59682 -76004 59734 -74866
rect 60036 -76012 60038 -74874
rect 60038 -76012 60092 -74874
rect 60386 -76010 60390 -74872
rect 60390 -76010 60442 -74872
rect 60748 -76006 60752 -74868
rect 60752 -76006 60804 -74868
rect 61102 -76010 61106 -74872
rect 61106 -76010 61158 -74872
rect 61460 -76004 61462 -74866
rect 61462 -76004 61516 -74866
rect 61810 -76010 61812 -74872
rect 61812 -76010 61866 -74872
rect 62172 -76012 62226 -74876
rect 62226 -76012 62228 -74876
rect 62172 -76014 62228 -76012
rect 62528 -76010 62530 -74872
rect 62530 -76010 62584 -74872
rect 62878 -76012 62882 -74876
rect 62882 -76012 62934 -74876
rect 62878 -76014 62934 -76012
rect 63238 -76006 63240 -74874
rect 63240 -76006 63294 -74874
rect 63238 -76012 63294 -76006
rect 63598 -76008 63650 -74876
rect 63650 -76008 63654 -74876
rect 63598 -76014 63654 -76008
rect 63950 -76006 63952 -74870
rect 63952 -76006 64006 -74870
rect 63950 -76008 64006 -76006
rect 64304 -76008 64306 -74870
rect 64306 -76008 64360 -74870
rect 56478 -78390 56480 -77252
rect 56480 -78390 56534 -77252
rect 56842 -78384 56896 -77246
rect 56896 -78384 56898 -77246
rect 57186 -78396 57192 -77258
rect 57192 -78396 57242 -77258
rect 57546 -78390 57548 -77252
rect 57548 -78390 57602 -77252
rect 57906 -78396 57960 -77258
rect 57960 -78396 57962 -77258
rect 58264 -78398 58266 -77260
rect 58266 -78398 58320 -77260
rect 58618 -77252 58674 -77250
rect 58618 -78388 58620 -77252
rect 58620 -78388 58674 -77252
rect 58970 -78392 58976 -77254
rect 58976 -78392 59026 -77254
rect 59332 -78388 59334 -77250
rect 59334 -78388 59388 -77250
rect 59684 -78392 59688 -77254
rect 59688 -78392 59740 -77254
rect 60042 -78400 60044 -77262
rect 60044 -78400 60098 -77262
rect 60392 -78398 60396 -77260
rect 60396 -78398 60448 -77260
rect 60754 -78394 60758 -77256
rect 60758 -78394 60810 -77256
rect 61108 -78398 61112 -77260
rect 61112 -78398 61164 -77260
rect 61466 -78392 61468 -77254
rect 61468 -78392 61522 -77254
rect 61816 -78398 61818 -77260
rect 61818 -78398 61872 -77260
rect 62178 -78400 62232 -77264
rect 62232 -78400 62234 -77264
rect 62178 -78402 62234 -78400
rect 62534 -78398 62536 -77260
rect 62536 -78398 62590 -77260
rect 62884 -78400 62888 -77264
rect 62888 -78400 62940 -77264
rect 62884 -78402 62940 -78400
rect 63244 -78394 63246 -77262
rect 63246 -78394 63300 -77262
rect 63244 -78400 63300 -78394
rect 63604 -78396 63656 -77264
rect 63656 -78396 63660 -77264
rect 63604 -78402 63660 -78396
rect 63956 -78394 63958 -77258
rect 63958 -78394 64012 -77258
rect 63956 -78396 64012 -78394
rect 64310 -78396 64312 -77258
rect 64312 -78396 64366 -77258
rect 56462 -79852 56464 -78714
rect 56464 -79852 56518 -78714
rect 56826 -79846 56880 -78708
rect 56880 -79846 56882 -78708
rect 57170 -79858 57176 -78720
rect 57176 -79858 57226 -78720
rect 57530 -79852 57532 -78714
rect 57532 -79852 57586 -78714
rect 57890 -79858 57944 -78720
rect 57944 -79858 57946 -78720
rect 58248 -79860 58250 -78722
rect 58250 -79860 58304 -78722
rect 58602 -78714 58658 -78712
rect 58602 -79850 58604 -78714
rect 58604 -79850 58658 -78714
rect 58954 -79854 58960 -78716
rect 58960 -79854 59010 -78716
rect 59316 -79850 59318 -78712
rect 59318 -79850 59372 -78712
rect 59668 -79854 59672 -78716
rect 59672 -79854 59724 -78716
rect 60026 -79862 60028 -78724
rect 60028 -79862 60082 -78724
rect 60376 -79860 60380 -78722
rect 60380 -79860 60432 -78722
rect 60738 -79856 60742 -78718
rect 60742 -79856 60794 -78718
rect 61092 -79860 61096 -78722
rect 61096 -79860 61148 -78722
rect 61450 -79854 61452 -78716
rect 61452 -79854 61506 -78716
rect 61800 -79860 61802 -78722
rect 61802 -79860 61856 -78722
rect 62162 -79862 62216 -78726
rect 62216 -79862 62218 -78726
rect 62162 -79864 62218 -79862
rect 62518 -79860 62520 -78722
rect 62520 -79860 62574 -78722
rect 62868 -79862 62872 -78726
rect 62872 -79862 62924 -78726
rect 62868 -79864 62924 -79862
rect 63228 -79856 63230 -78724
rect 63230 -79856 63284 -78724
rect 63228 -79862 63284 -79856
rect 63588 -79858 63640 -78726
rect 63640 -79858 63644 -78726
rect 63588 -79864 63644 -79858
rect 63940 -79856 63942 -78720
rect 63942 -79856 63996 -78720
rect 63940 -79858 63996 -79856
rect 64294 -79858 64296 -78720
rect 64296 -79858 64350 -78720
rect 56488 -82356 56490 -81218
rect 56490 -82356 56544 -81218
rect 56852 -82350 56906 -81212
rect 56906 -82350 56908 -81212
rect 57196 -82362 57202 -81224
rect 57202 -82362 57252 -81224
rect 57556 -82356 57558 -81218
rect 57558 -82356 57612 -81218
rect 57916 -82362 57970 -81224
rect 57970 -82362 57972 -81224
rect 58274 -82364 58276 -81226
rect 58276 -82364 58330 -81226
rect 58628 -81218 58684 -81216
rect 58628 -82354 58630 -81218
rect 58630 -82354 58684 -81218
rect 58980 -82358 58986 -81220
rect 58986 -82358 59036 -81220
rect 59342 -82354 59344 -81216
rect 59344 -82354 59398 -81216
rect 59694 -82358 59698 -81220
rect 59698 -82358 59750 -81220
rect 60052 -82366 60054 -81228
rect 60054 -82366 60108 -81228
rect 60402 -82364 60406 -81226
rect 60406 -82364 60458 -81226
rect 60764 -82360 60768 -81222
rect 60768 -82360 60820 -81222
rect 61118 -82364 61122 -81226
rect 61122 -82364 61174 -81226
rect 61476 -82358 61478 -81220
rect 61478 -82358 61532 -81220
rect 61826 -82364 61828 -81226
rect 61828 -82364 61882 -81226
rect 62188 -82366 62242 -81230
rect 62242 -82366 62244 -81230
rect 62188 -82368 62244 -82366
rect 62544 -82364 62546 -81226
rect 62546 -82364 62600 -81226
rect 62894 -82366 62898 -81230
rect 62898 -82366 62950 -81230
rect 62894 -82368 62950 -82366
rect 63254 -82360 63256 -81228
rect 63256 -82360 63310 -81228
rect 63254 -82366 63310 -82360
rect 63614 -82362 63666 -81230
rect 63666 -82362 63670 -81230
rect 63614 -82368 63670 -82362
rect 63966 -82360 63968 -81224
rect 63968 -82360 64022 -81224
rect 63966 -82362 64022 -82360
rect 64320 -82362 64322 -81224
rect 64322 -82362 64376 -81224
rect 56472 -83818 56474 -82680
rect 56474 -83818 56528 -82680
rect 56836 -83812 56890 -82674
rect 56890 -83812 56892 -82674
rect 57180 -83824 57186 -82686
rect 57186 -83824 57236 -82686
rect 57540 -83818 57542 -82680
rect 57542 -83818 57596 -82680
rect 57900 -83824 57954 -82686
rect 57954 -83824 57956 -82686
rect 58258 -83826 58260 -82688
rect 58260 -83826 58314 -82688
rect 58612 -82680 58668 -82678
rect 58612 -83816 58614 -82680
rect 58614 -83816 58668 -82680
rect 58964 -83820 58970 -82682
rect 58970 -83820 59020 -82682
rect 59326 -83816 59328 -82678
rect 59328 -83816 59382 -82678
rect 59678 -83820 59682 -82682
rect 59682 -83820 59734 -82682
rect 60036 -83828 60038 -82690
rect 60038 -83828 60092 -82690
rect 60386 -83826 60390 -82688
rect 60390 -83826 60442 -82688
rect 60748 -83822 60752 -82684
rect 60752 -83822 60804 -82684
rect 61102 -83826 61106 -82688
rect 61106 -83826 61158 -82688
rect 61460 -83820 61462 -82682
rect 61462 -83820 61516 -82682
rect 61810 -83826 61812 -82688
rect 61812 -83826 61866 -82688
rect 62172 -83828 62226 -82692
rect 62226 -83828 62228 -82692
rect 62172 -83830 62228 -83828
rect 62528 -83826 62530 -82688
rect 62530 -83826 62584 -82688
rect 62878 -83828 62882 -82692
rect 62882 -83828 62934 -82692
rect 62878 -83830 62934 -83828
rect 63238 -83822 63240 -82690
rect 63240 -83822 63294 -82690
rect 63238 -83828 63294 -83822
rect 63598 -83824 63650 -82692
rect 63650 -83824 63654 -82692
rect 63598 -83830 63654 -83824
rect 63950 -83822 63952 -82686
rect 63952 -83822 64006 -82686
rect 63950 -83824 64006 -83822
rect 64304 -83824 64306 -82686
rect 64306 -83824 64360 -82686
rect 56460 -86176 56462 -85038
rect 56462 -86176 56516 -85038
rect 56824 -86170 56878 -85032
rect 56878 -86170 56880 -85032
rect 57168 -86182 57174 -85044
rect 57174 -86182 57224 -85044
rect 57528 -86176 57530 -85038
rect 57530 -86176 57584 -85038
rect 57888 -86182 57942 -85044
rect 57942 -86182 57944 -85044
rect 58246 -86184 58248 -85046
rect 58248 -86184 58302 -85046
rect 58600 -85038 58656 -85036
rect 58600 -86174 58602 -85038
rect 58602 -86174 58656 -85038
rect 58952 -86178 58958 -85040
rect 58958 -86178 59008 -85040
rect 59314 -86174 59316 -85036
rect 59316 -86174 59370 -85036
rect 59666 -86178 59670 -85040
rect 59670 -86178 59722 -85040
rect 60024 -86186 60026 -85048
rect 60026 -86186 60080 -85048
rect 60374 -86184 60378 -85046
rect 60378 -86184 60430 -85046
rect 60736 -86180 60740 -85042
rect 60740 -86180 60792 -85042
rect 61090 -86184 61094 -85046
rect 61094 -86184 61146 -85046
rect 61448 -86178 61450 -85040
rect 61450 -86178 61504 -85040
rect 61798 -86184 61800 -85046
rect 61800 -86184 61854 -85046
rect 62160 -86186 62214 -85050
rect 62214 -86186 62216 -85050
rect 62160 -86188 62216 -86186
rect 62516 -86184 62518 -85046
rect 62518 -86184 62572 -85046
rect 62866 -86186 62870 -85050
rect 62870 -86186 62922 -85050
rect 62866 -86188 62922 -86186
rect 63226 -86180 63228 -85048
rect 63228 -86180 63282 -85048
rect 63226 -86186 63282 -86180
rect 63586 -86182 63638 -85050
rect 63638 -86182 63642 -85050
rect 63586 -86188 63642 -86182
rect 63938 -86180 63940 -85044
rect 63940 -86180 63994 -85044
rect 63938 -86182 63994 -86180
rect 64292 -86182 64294 -85044
rect 64294 -86182 64348 -85044
rect 56444 -87638 56446 -86500
rect 56446 -87638 56500 -86500
rect 56808 -87632 56862 -86494
rect 56862 -87632 56864 -86494
rect 57152 -87644 57158 -86506
rect 57158 -87644 57208 -86506
rect 57512 -87638 57514 -86500
rect 57514 -87638 57568 -86500
rect 57872 -87644 57926 -86506
rect 57926 -87644 57928 -86506
rect 58230 -87646 58232 -86508
rect 58232 -87646 58286 -86508
rect 58584 -86500 58640 -86498
rect 58584 -87636 58586 -86500
rect 58586 -87636 58640 -86500
rect 58936 -87640 58942 -86502
rect 58942 -87640 58992 -86502
rect 59298 -87636 59300 -86498
rect 59300 -87636 59354 -86498
rect 59650 -87640 59654 -86502
rect 59654 -87640 59706 -86502
rect 60008 -87648 60010 -86510
rect 60010 -87648 60064 -86510
rect 60358 -87646 60362 -86508
rect 60362 -87646 60414 -86508
rect 60720 -87642 60724 -86504
rect 60724 -87642 60776 -86504
rect 61074 -87646 61078 -86508
rect 61078 -87646 61130 -86508
rect 61432 -87640 61434 -86502
rect 61434 -87640 61488 -86502
rect 61782 -87646 61784 -86508
rect 61784 -87646 61838 -86508
rect 62144 -87648 62198 -86512
rect 62198 -87648 62200 -86512
rect 62144 -87650 62200 -87648
rect 62500 -87646 62502 -86508
rect 62502 -87646 62556 -86508
rect 62850 -87648 62854 -86512
rect 62854 -87648 62906 -86512
rect 62850 -87650 62906 -87648
rect 63210 -87642 63212 -86510
rect 63212 -87642 63266 -86510
rect 63210 -87648 63266 -87642
rect 63570 -87644 63622 -86512
rect 63622 -87644 63626 -86512
rect 63570 -87650 63626 -87644
rect 63922 -87642 63924 -86506
rect 63924 -87642 63978 -86506
rect 63922 -87644 63978 -87642
rect 64276 -87644 64278 -86506
rect 64278 -87644 64332 -86506
rect 66316 -87788 66318 -87634
rect 66318 -87788 66372 -87634
rect 66674 -87788 66676 -87634
rect 66676 -87788 66730 -87634
rect 67028 -87786 67030 -87632
rect 67030 -87786 67084 -87632
rect 66324 -88214 66326 -88060
rect 66326 -88214 66380 -88060
rect 66702 -88216 66740 -88070
rect 66740 -88216 66758 -88070
rect 66702 -88224 66758 -88216
rect 67038 -88216 67040 -88062
rect 67040 -88216 67094 -88062
rect 66318 -88620 66320 -88466
rect 66320 -88620 66374 -88466
rect 66674 -88626 66676 -88472
rect 66676 -88626 66730 -88472
rect 67032 -88622 67034 -88468
rect 67034 -88622 67088 -88468
rect 66318 -89034 66320 -88880
rect 66320 -89034 66372 -88880
rect 66372 -89034 66374 -88880
rect 66670 -89034 66672 -88880
rect 66672 -89034 66724 -88880
rect 66724 -89034 66726 -88880
rect 67032 -89034 67034 -88880
rect 67034 -89034 67086 -88880
rect 67086 -89034 67088 -88880
rect 68260 -87882 68318 -87872
rect 68260 -89018 68312 -87882
rect 68312 -89018 68318 -87882
rect 68260 -89024 68318 -89018
rect 68440 -87876 68498 -87868
rect 68440 -89012 68442 -87876
rect 68442 -89012 68494 -87876
rect 68494 -89012 68498 -87876
rect 68440 -89020 68498 -89012
rect 68628 -87884 68686 -87868
rect 68628 -89020 68680 -87884
rect 68680 -89020 68686 -87884
rect 68802 -87890 68860 -87874
rect 68802 -89026 68854 -87890
rect 68854 -89026 68860 -87890
rect 68978 -87890 69036 -87872
rect 68978 -89024 68980 -87890
rect 68980 -89024 69032 -87890
rect 69032 -89024 69036 -87890
rect 69160 -87890 69218 -87874
rect 69160 -89026 69212 -87890
rect 69212 -89026 69218 -87890
rect 69338 -87890 69396 -87874
rect 69338 -89026 69388 -87890
rect 69388 -89026 69396 -87890
rect 69512 -87886 69570 -87872
rect 69512 -89022 69514 -87886
rect 69514 -89022 69566 -87886
rect 69566 -89022 69570 -87886
rect 69512 -89024 69570 -89022
rect 69692 -87888 69750 -87872
rect 69692 -89024 69694 -87888
rect 69694 -89024 69746 -87888
rect 69746 -89024 69750 -87888
rect 69866 -87886 69924 -87874
rect 69866 -89022 69868 -87886
rect 69868 -89022 69920 -87886
rect 69920 -89022 69924 -87886
rect 69866 -89026 69924 -89022
rect 70048 -87890 70106 -87878
rect 70048 -89026 70100 -87890
rect 70100 -89026 70106 -87890
rect 70048 -89030 70106 -89026
rect 70222 -87888 70280 -87880
rect 70222 -89024 70224 -87888
rect 70224 -89024 70276 -87888
rect 70276 -89024 70280 -87888
rect 70222 -89032 70280 -89024
rect 70400 -87888 70458 -87872
rect 70400 -89024 70404 -87888
rect 70404 -89024 70456 -87888
rect 70456 -89024 70458 -87888
rect 70582 -87890 70640 -87878
rect 70582 -89026 70634 -87890
rect 70634 -89026 70640 -87890
rect 70582 -89030 70640 -89026
rect 70756 -87892 70814 -87878
rect 70756 -89028 70760 -87892
rect 70760 -89028 70812 -87892
rect 70812 -89028 70814 -87892
rect 70756 -89030 70814 -89028
rect 70936 -87890 70994 -87876
rect 70936 -89026 70988 -87890
rect 70988 -89026 70994 -87890
rect 70936 -89028 70994 -89026
rect 71118 -87892 71176 -87876
rect 71118 -89028 71166 -87892
rect 71166 -89028 71176 -87892
rect 71292 -87890 71350 -87882
rect 71292 -89026 71294 -87890
rect 71294 -89026 71346 -87890
rect 71346 -89026 71350 -87890
rect 71292 -89034 71350 -89026
rect 71472 -87890 71530 -87880
rect 71472 -89026 71524 -87890
rect 71524 -89026 71530 -87890
rect 71472 -89032 71530 -89026
rect 71646 -87892 71704 -87880
rect 71646 -89028 71648 -87892
rect 71648 -89028 71700 -87892
rect 71700 -89028 71704 -87892
rect 71646 -89032 71704 -89028
rect 71824 -87890 71882 -87876
rect 71824 -89026 71826 -87890
rect 71826 -89026 71878 -87890
rect 71878 -89026 71882 -87890
rect 71824 -89028 71882 -89026
rect 74156 -87880 74214 -87870
rect 74156 -89016 74208 -87880
rect 74208 -89016 74214 -87880
rect 74156 -89022 74214 -89016
rect 74336 -87874 74394 -87866
rect 74336 -89010 74338 -87874
rect 74338 -89010 74390 -87874
rect 74390 -89010 74394 -87874
rect 74336 -89018 74394 -89010
rect 74524 -87882 74582 -87866
rect 74524 -89018 74576 -87882
rect 74576 -89018 74582 -87882
rect 74698 -87888 74756 -87872
rect 74698 -89024 74750 -87888
rect 74750 -89024 74756 -87888
rect 74874 -87888 74932 -87870
rect 74874 -89022 74876 -87888
rect 74876 -89022 74928 -87888
rect 74928 -89022 74932 -87888
rect 75056 -87888 75114 -87872
rect 75056 -89024 75108 -87888
rect 75108 -89024 75114 -87888
rect 75234 -87888 75292 -87872
rect 75234 -89024 75284 -87888
rect 75284 -89024 75292 -87888
rect 75408 -87884 75466 -87870
rect 75408 -89020 75410 -87884
rect 75410 -89020 75462 -87884
rect 75462 -89020 75466 -87884
rect 75408 -89022 75466 -89020
rect 75588 -87886 75646 -87870
rect 75588 -89022 75590 -87886
rect 75590 -89022 75642 -87886
rect 75642 -89022 75646 -87886
rect 75762 -87884 75820 -87872
rect 75762 -89020 75764 -87884
rect 75764 -89020 75816 -87884
rect 75816 -89020 75820 -87884
rect 75762 -89024 75820 -89020
rect 75944 -87888 76002 -87876
rect 75944 -89024 75996 -87888
rect 75996 -89024 76002 -87888
rect 75944 -89028 76002 -89024
rect 76118 -87886 76176 -87878
rect 76118 -89022 76120 -87886
rect 76120 -89022 76172 -87886
rect 76172 -89022 76176 -87886
rect 76118 -89030 76176 -89022
rect 76296 -87886 76354 -87870
rect 76296 -89022 76300 -87886
rect 76300 -89022 76352 -87886
rect 76352 -89022 76354 -87886
rect 76478 -87888 76536 -87876
rect 76478 -89024 76530 -87888
rect 76530 -89024 76536 -87888
rect 76478 -89028 76536 -89024
rect 76652 -87890 76710 -87876
rect 76652 -89026 76656 -87890
rect 76656 -89026 76708 -87890
rect 76708 -89026 76710 -87890
rect 76652 -89028 76710 -89026
rect 76832 -87888 76890 -87874
rect 76832 -89024 76884 -87888
rect 76884 -89024 76890 -87888
rect 76832 -89026 76890 -89024
rect 77014 -87890 77072 -87874
rect 77014 -89026 77062 -87890
rect 77062 -89026 77072 -87890
rect 77188 -87888 77246 -87880
rect 77188 -89024 77190 -87888
rect 77190 -89024 77242 -87888
rect 77242 -89024 77246 -87888
rect 77188 -89032 77246 -89024
rect 77368 -87888 77426 -87878
rect 77368 -89024 77420 -87888
rect 77420 -89024 77426 -87888
rect 77368 -89030 77426 -89024
rect 77542 -87890 77600 -87878
rect 77542 -89026 77544 -87890
rect 77544 -89026 77596 -87890
rect 77596 -89026 77600 -87890
rect 77542 -89030 77600 -89026
rect 77720 -87888 77778 -87874
rect 77720 -89024 77722 -87888
rect 77722 -89024 77774 -87888
rect 77774 -89024 77778 -87888
rect 77720 -89026 77778 -89024
rect 80270 -87874 80328 -87864
rect 80270 -89010 80322 -87874
rect 80322 -89010 80328 -87874
rect 80270 -89016 80328 -89010
rect 80450 -87868 80508 -87860
rect 80450 -89004 80452 -87868
rect 80452 -89004 80504 -87868
rect 80504 -89004 80508 -87868
rect 80450 -89012 80508 -89004
rect 80638 -87876 80696 -87860
rect 80638 -89012 80690 -87876
rect 80690 -89012 80696 -87876
rect 80812 -87882 80870 -87866
rect 80812 -89018 80864 -87882
rect 80864 -89018 80870 -87882
rect 80988 -87882 81046 -87864
rect 80988 -89016 80990 -87882
rect 80990 -89016 81042 -87882
rect 81042 -89016 81046 -87882
rect 81170 -87882 81228 -87866
rect 81170 -89018 81222 -87882
rect 81222 -89018 81228 -87882
rect 81348 -87882 81406 -87866
rect 81348 -89018 81398 -87882
rect 81398 -89018 81406 -87882
rect 81522 -87878 81580 -87864
rect 81522 -89014 81524 -87878
rect 81524 -89014 81576 -87878
rect 81576 -89014 81580 -87878
rect 81522 -89016 81580 -89014
rect 81702 -87880 81760 -87864
rect 81702 -89016 81704 -87880
rect 81704 -89016 81756 -87880
rect 81756 -89016 81760 -87880
rect 81876 -87878 81934 -87866
rect 81876 -89014 81878 -87878
rect 81878 -89014 81930 -87878
rect 81930 -89014 81934 -87878
rect 81876 -89018 81934 -89014
rect 82058 -87882 82116 -87870
rect 82058 -89018 82110 -87882
rect 82110 -89018 82116 -87882
rect 82058 -89022 82116 -89018
rect 82232 -87880 82290 -87872
rect 82232 -89016 82234 -87880
rect 82234 -89016 82286 -87880
rect 82286 -89016 82290 -87880
rect 82232 -89024 82290 -89016
rect 82410 -87880 82468 -87864
rect 82410 -89016 82414 -87880
rect 82414 -89016 82466 -87880
rect 82466 -89016 82468 -87880
rect 82592 -87882 82650 -87870
rect 82592 -89018 82644 -87882
rect 82644 -89018 82650 -87882
rect 82592 -89022 82650 -89018
rect 82766 -87884 82824 -87870
rect 82766 -89020 82770 -87884
rect 82770 -89020 82822 -87884
rect 82822 -89020 82824 -87884
rect 82766 -89022 82824 -89020
rect 82946 -87882 83004 -87868
rect 82946 -89018 82998 -87882
rect 82998 -89018 83004 -87882
rect 82946 -89020 83004 -89018
rect 83128 -87884 83186 -87868
rect 83128 -89020 83176 -87884
rect 83176 -89020 83186 -87884
rect 83302 -87882 83360 -87874
rect 83302 -89018 83304 -87882
rect 83304 -89018 83356 -87882
rect 83356 -89018 83360 -87882
rect 83302 -89026 83360 -89018
rect 83482 -87882 83540 -87872
rect 83482 -89018 83534 -87882
rect 83534 -89018 83540 -87882
rect 83482 -89024 83540 -89018
rect 83656 -87884 83714 -87872
rect 83656 -89020 83658 -87884
rect 83658 -89020 83710 -87884
rect 83710 -89020 83714 -87884
rect 83656 -89024 83714 -89020
rect 83834 -87882 83892 -87868
rect 83834 -89018 83836 -87882
rect 83836 -89018 83888 -87882
rect 83888 -89018 83892 -87882
rect 83834 -89020 83892 -89018
rect 56542 -90472 56548 -89338
rect 56548 -90472 56600 -89338
rect 56600 -90472 56602 -89338
rect 56900 -90470 56906 -89336
rect 56906 -90470 56958 -89336
rect 56958 -90470 56960 -89336
rect 57254 -90476 57260 -89342
rect 57260 -90476 57312 -89342
rect 57312 -90476 57314 -89342
rect 57608 -90482 57614 -89348
rect 57614 -90482 57666 -89348
rect 57666 -90482 57668 -89348
rect 57964 -90478 57974 -89344
rect 57974 -90478 58024 -89344
rect 58322 -90474 58328 -89340
rect 58328 -90474 58380 -89340
rect 58380 -90474 58382 -89340
rect 58682 -90468 58686 -89334
rect 58686 -90468 58738 -89334
rect 58738 -90468 58742 -89334
rect 59028 -90480 59038 -89346
rect 59038 -90480 59088 -89346
rect 59388 -90472 59396 -89338
rect 59396 -90472 59448 -89338
rect 59746 -90464 59752 -89330
rect 59752 -90464 59804 -89330
rect 59804 -90464 59806 -89330
rect 60974 -90474 60980 -89340
rect 60980 -90474 61032 -89340
rect 61032 -90474 61034 -89340
rect 61322 -90476 61330 -89342
rect 61330 -90476 61382 -89342
rect 61680 -90468 61690 -89334
rect 61690 -90468 61740 -89334
rect 62042 -90478 62094 -89344
rect 62094 -90478 62102 -89344
rect 62396 -90482 62398 -89348
rect 62398 -90482 62450 -89348
rect 62450 -90482 62456 -89348
rect 62752 -90482 62756 -89348
rect 62756 -90482 62808 -89348
rect 62808 -90482 62812 -89348
rect 63106 -90474 63112 -89340
rect 63112 -90474 63164 -89340
rect 63164 -90474 63166 -89340
rect 63466 -90486 63468 -89352
rect 63468 -90486 63520 -89352
rect 63520 -90486 63526 -89352
rect 63826 -90478 63878 -89344
rect 63878 -90478 63886 -89344
rect 64182 -90482 64184 -89348
rect 64184 -90482 64236 -89348
rect 64236 -90482 64242 -89348
rect 68268 -89308 68326 -89300
rect 68268 -90444 68320 -89308
rect 68320 -90444 68326 -89308
rect 68268 -90452 68326 -90444
rect 68444 -89308 68502 -89294
rect 68444 -90444 68446 -89308
rect 68446 -90444 68498 -89308
rect 68498 -90444 68502 -89308
rect 68444 -90446 68502 -90444
rect 68622 -89306 68680 -89290
rect 68622 -90442 68672 -89306
rect 68672 -90442 68680 -89306
rect 68800 -89310 68858 -89296
rect 68800 -90446 68802 -89310
rect 68802 -90446 68854 -89310
rect 68854 -90446 68858 -89310
rect 68800 -90448 68858 -90446
rect 68980 -89308 69038 -89298
rect 68980 -90444 69032 -89308
rect 69032 -90444 69038 -89308
rect 68980 -90450 69038 -90444
rect 69156 -89306 69214 -89294
rect 69156 -90442 69208 -89306
rect 69208 -90442 69214 -89306
rect 69156 -90446 69214 -90442
rect 69332 -89310 69390 -89298
rect 69332 -90446 69334 -89310
rect 69334 -90446 69386 -89310
rect 69386 -90446 69390 -89310
rect 69332 -90450 69390 -90446
rect 69508 -89308 69566 -89292
rect 69508 -90444 69512 -89308
rect 69512 -90444 69564 -89308
rect 69564 -90444 69566 -89308
rect 69688 -89306 69746 -89294
rect 69688 -90442 69690 -89306
rect 69690 -90442 69742 -89306
rect 69742 -90442 69746 -89306
rect 69688 -90446 69746 -90442
rect 69864 -89310 69922 -89298
rect 69864 -90446 69866 -89310
rect 69866 -90446 69918 -89310
rect 69918 -90446 69922 -89310
rect 69864 -90450 69922 -90446
rect 70044 -89308 70102 -89294
rect 70044 -90444 70046 -89308
rect 70046 -90444 70098 -89308
rect 70098 -90444 70102 -89308
rect 70044 -90446 70102 -90444
rect 70226 -89308 70284 -89292
rect 70226 -90444 70278 -89308
rect 70278 -90444 70284 -89308
rect 70406 -89308 70464 -89294
rect 70406 -90444 70458 -89308
rect 70458 -90444 70464 -89308
rect 70406 -90446 70464 -90444
rect 70578 -89308 70636 -89294
rect 70578 -90444 70580 -89308
rect 70580 -90444 70632 -89308
rect 70632 -90444 70636 -89308
rect 70578 -90446 70636 -90444
rect 70756 -89306 70814 -89294
rect 70756 -90442 70758 -89306
rect 70758 -90442 70810 -89306
rect 70810 -90442 70814 -89306
rect 70756 -90446 70814 -90442
rect 70934 -89306 70992 -89294
rect 70934 -90442 70986 -89306
rect 70986 -90442 70992 -89306
rect 70934 -90446 70992 -90442
rect 71112 -89306 71170 -89288
rect 71112 -90440 71114 -89306
rect 71114 -90440 71166 -89306
rect 71166 -90440 71170 -89306
rect 71294 -89312 71352 -89298
rect 71294 -90448 71344 -89312
rect 71344 -90448 71352 -89312
rect 71294 -90450 71352 -90448
rect 71472 -89308 71530 -89300
rect 71472 -90444 71524 -89308
rect 71524 -90444 71530 -89308
rect 71472 -90452 71530 -90444
rect 71646 -89310 71704 -89294
rect 71646 -90446 71648 -89310
rect 71648 -90446 71700 -89310
rect 71700 -90446 71704 -89310
rect 71826 -89310 71884 -89298
rect 71826 -90446 71878 -89310
rect 71878 -90446 71884 -89310
rect 71826 -90450 71884 -90446
rect 74164 -89306 74222 -89298
rect 74164 -90442 74216 -89306
rect 74216 -90442 74222 -89306
rect 74164 -90450 74222 -90442
rect 74340 -89306 74398 -89292
rect 74340 -90442 74342 -89306
rect 74342 -90442 74394 -89306
rect 74394 -90442 74398 -89306
rect 74340 -90444 74398 -90442
rect 74518 -89304 74576 -89288
rect 74518 -90440 74568 -89304
rect 74568 -90440 74576 -89304
rect 74696 -89308 74754 -89294
rect 74696 -90444 74698 -89308
rect 74698 -90444 74750 -89308
rect 74750 -90444 74754 -89308
rect 74696 -90446 74754 -90444
rect 74876 -89306 74934 -89296
rect 74876 -90442 74928 -89306
rect 74928 -90442 74934 -89306
rect 74876 -90448 74934 -90442
rect 75052 -89304 75110 -89292
rect 75052 -90440 75104 -89304
rect 75104 -90440 75110 -89304
rect 75052 -90444 75110 -90440
rect 75228 -89308 75286 -89296
rect 75228 -90444 75230 -89308
rect 75230 -90444 75282 -89308
rect 75282 -90444 75286 -89308
rect 75228 -90448 75286 -90444
rect 75404 -89306 75462 -89290
rect 75404 -90442 75408 -89306
rect 75408 -90442 75460 -89306
rect 75460 -90442 75462 -89306
rect 75584 -89304 75642 -89292
rect 75584 -90440 75586 -89304
rect 75586 -90440 75638 -89304
rect 75638 -90440 75642 -89304
rect 75584 -90444 75642 -90440
rect 75760 -89308 75818 -89296
rect 75760 -90444 75762 -89308
rect 75762 -90444 75814 -89308
rect 75814 -90444 75818 -89308
rect 75760 -90448 75818 -90444
rect 75940 -89306 75998 -89292
rect 75940 -90442 75942 -89306
rect 75942 -90442 75994 -89306
rect 75994 -90442 75998 -89306
rect 75940 -90444 75998 -90442
rect 76122 -89306 76180 -89290
rect 76122 -90442 76174 -89306
rect 76174 -90442 76180 -89306
rect 76302 -89306 76360 -89292
rect 76302 -90442 76354 -89306
rect 76354 -90442 76360 -89306
rect 76302 -90444 76360 -90442
rect 76474 -89306 76532 -89292
rect 76474 -90442 76476 -89306
rect 76476 -90442 76528 -89306
rect 76528 -90442 76532 -89306
rect 76474 -90444 76532 -90442
rect 76652 -89304 76710 -89292
rect 76652 -90440 76654 -89304
rect 76654 -90440 76706 -89304
rect 76706 -90440 76710 -89304
rect 76652 -90444 76710 -90440
rect 76830 -89304 76888 -89292
rect 76830 -90440 76882 -89304
rect 76882 -90440 76888 -89304
rect 76830 -90444 76888 -90440
rect 77008 -89304 77066 -89286
rect 77008 -90438 77010 -89304
rect 77010 -90438 77062 -89304
rect 77062 -90438 77066 -89304
rect 77190 -89310 77248 -89296
rect 77190 -90446 77240 -89310
rect 77240 -90446 77248 -89310
rect 77190 -90448 77248 -90446
rect 77368 -89306 77426 -89298
rect 77368 -90442 77420 -89306
rect 77420 -90442 77426 -89306
rect 77368 -90450 77426 -90442
rect 77542 -89308 77600 -89292
rect 77542 -90444 77544 -89308
rect 77544 -90444 77596 -89308
rect 77596 -90444 77600 -89308
rect 77722 -89308 77780 -89296
rect 77722 -90444 77774 -89308
rect 77774 -90444 77780 -89308
rect 77722 -90448 77780 -90444
rect 80278 -89300 80336 -89292
rect 80278 -90436 80330 -89300
rect 80330 -90436 80336 -89300
rect 80278 -90444 80336 -90436
rect 80454 -89300 80512 -89286
rect 80454 -90436 80456 -89300
rect 80456 -90436 80508 -89300
rect 80508 -90436 80512 -89300
rect 80454 -90438 80512 -90436
rect 80632 -89298 80690 -89282
rect 80632 -90434 80682 -89298
rect 80682 -90434 80690 -89298
rect 80810 -89302 80868 -89288
rect 80810 -90438 80812 -89302
rect 80812 -90438 80864 -89302
rect 80864 -90438 80868 -89302
rect 80810 -90440 80868 -90438
rect 80990 -89300 81048 -89290
rect 80990 -90436 81042 -89300
rect 81042 -90436 81048 -89300
rect 80990 -90442 81048 -90436
rect 81166 -89298 81224 -89286
rect 81166 -90434 81218 -89298
rect 81218 -90434 81224 -89298
rect 81166 -90438 81224 -90434
rect 81342 -89302 81400 -89290
rect 81342 -90438 81344 -89302
rect 81344 -90438 81396 -89302
rect 81396 -90438 81400 -89302
rect 81342 -90442 81400 -90438
rect 81518 -89300 81576 -89284
rect 81518 -90436 81522 -89300
rect 81522 -90436 81574 -89300
rect 81574 -90436 81576 -89300
rect 81698 -89298 81756 -89286
rect 81698 -90434 81700 -89298
rect 81700 -90434 81752 -89298
rect 81752 -90434 81756 -89298
rect 81698 -90438 81756 -90434
rect 81874 -89302 81932 -89290
rect 81874 -90438 81876 -89302
rect 81876 -90438 81928 -89302
rect 81928 -90438 81932 -89302
rect 81874 -90442 81932 -90438
rect 82054 -89300 82112 -89286
rect 82054 -90436 82056 -89300
rect 82056 -90436 82108 -89300
rect 82108 -90436 82112 -89300
rect 82054 -90438 82112 -90436
rect 82236 -89300 82294 -89284
rect 82236 -90436 82288 -89300
rect 82288 -90436 82294 -89300
rect 82416 -89300 82474 -89286
rect 82416 -90436 82468 -89300
rect 82468 -90436 82474 -89300
rect 82416 -90438 82474 -90436
rect 82588 -89300 82646 -89286
rect 82588 -90436 82590 -89300
rect 82590 -90436 82642 -89300
rect 82642 -90436 82646 -89300
rect 82588 -90438 82646 -90436
rect 82766 -89298 82824 -89286
rect 82766 -90434 82768 -89298
rect 82768 -90434 82820 -89298
rect 82820 -90434 82824 -89298
rect 82766 -90438 82824 -90434
rect 82944 -89298 83002 -89286
rect 82944 -90434 82996 -89298
rect 82996 -90434 83002 -89298
rect 82944 -90438 83002 -90434
rect 83122 -89298 83180 -89280
rect 83122 -90432 83124 -89298
rect 83124 -90432 83176 -89298
rect 83176 -90432 83180 -89298
rect 83304 -89304 83362 -89290
rect 83304 -90440 83354 -89304
rect 83354 -90440 83362 -89304
rect 83304 -90442 83362 -90440
rect 83482 -89300 83540 -89292
rect 83482 -90436 83534 -89300
rect 83534 -90436 83540 -89300
rect 83482 -90444 83540 -90436
rect 83656 -89302 83714 -89286
rect 83656 -90438 83658 -89302
rect 83658 -90438 83710 -89302
rect 83710 -90438 83714 -89302
rect 83836 -89302 83894 -89290
rect 83836 -90438 83888 -89302
rect 83888 -90438 83894 -89302
rect 83836 -90442 83894 -90438
<< metal3 >>
rect 60928 -70129 61004 -70120
rect 60928 -70134 61026 -70129
rect 60928 -71284 60946 -70134
rect 61016 -71284 61026 -70134
rect 60928 -71289 61026 -71284
rect 61286 -70133 61362 -70114
rect 61286 -70138 61382 -70133
rect 61286 -71288 61302 -70138
rect 61372 -71288 61382 -70138
rect 60928 -72630 61004 -71289
rect 61286 -71293 61382 -71288
rect 61642 -70137 61718 -70116
rect 62004 -70125 62080 -70114
rect 61994 -70130 62084 -70125
rect 61642 -70142 61734 -70137
rect 61642 -71292 61654 -70142
rect 61724 -71292 61734 -70142
rect 61994 -71280 62004 -70130
rect 62074 -71280 62084 -70130
rect 61994 -71285 62084 -71280
rect 62348 -70139 62424 -70122
rect 62710 -70137 62786 -70114
rect 63070 -70125 63146 -70120
rect 63414 -70125 63490 -70120
rect 63780 -70123 63856 -70116
rect 64140 -70122 64230 -70119
rect 63070 -70130 63168 -70125
rect 62348 -70144 62446 -70139
rect 61286 -72630 61362 -71293
rect 61642 -71297 61734 -71292
rect 61642 -72630 61718 -71297
rect 62004 -72630 62080 -71285
rect 62348 -71294 62366 -70144
rect 62436 -71294 62446 -70144
rect 62348 -71299 62446 -71294
rect 62710 -70142 62806 -70137
rect 62710 -71292 62726 -70142
rect 62796 -71292 62806 -70142
rect 62710 -71297 62806 -71292
rect 63070 -71280 63088 -70130
rect 63158 -71280 63168 -70130
rect 63070 -71285 63168 -71280
rect 63414 -70130 63516 -70125
rect 63414 -71280 63436 -70130
rect 63506 -71280 63516 -70130
rect 63414 -71285 63516 -71280
rect 63780 -70128 63874 -70123
rect 63780 -71278 63794 -70128
rect 63864 -71278 63874 -70128
rect 63780 -71283 63874 -71278
rect 64134 -70124 64230 -70122
rect 64134 -71274 64150 -70124
rect 64220 -71274 64230 -70124
rect 68304 -71268 68314 -70086
rect 68390 -71268 68400 -70086
rect 68656 -71268 68666 -70086
rect 68742 -71268 68752 -70086
rect 69010 -71260 69020 -70078
rect 69096 -71260 69106 -70078
rect 69016 -71265 69098 -71260
rect 69366 -71262 69376 -70080
rect 69452 -71262 69462 -70080
rect 69718 -71262 69728 -70080
rect 69804 -71262 69814 -70080
rect 69368 -71264 69378 -71262
rect 69440 -71264 69450 -71262
rect 64134 -71279 64230 -71274
rect 68310 -71270 68320 -71268
rect 68382 -71270 68392 -71268
rect 68310 -71275 68392 -71270
rect 68660 -71271 68742 -71268
rect 69368 -71269 69450 -71264
rect 69722 -71267 69804 -71262
rect 70080 -71274 70090 -70092
rect 70166 -71274 70176 -70092
rect 70434 -71260 70444 -70078
rect 70520 -71260 70530 -70078
rect 70782 -71252 70792 -70070
rect 70868 -71252 70878 -70070
rect 70794 -71254 70804 -71252
rect 70866 -71254 70876 -71252
rect 70794 -71259 70876 -71254
rect 71140 -71260 71150 -70078
rect 71226 -71260 71236 -70078
rect 70442 -71263 70524 -71260
rect 71148 -71263 71230 -71260
rect 71496 -71262 71506 -70080
rect 71582 -71262 71592 -70080
rect 71858 -71260 71868 -70078
rect 71944 -71260 71954 -70078
rect 72212 -71260 72222 -70078
rect 72298 -71260 72308 -70078
rect 72574 -71256 72584 -70074
rect 72660 -71256 72670 -70074
rect 71502 -71263 71584 -71262
rect 71864 -71263 71946 -71260
rect 72218 -71262 72228 -71260
rect 72290 -71262 72300 -71260
rect 72218 -71267 72300 -71262
rect 72576 -71262 72586 -71256
rect 72648 -71262 72658 -71256
rect 72928 -71258 72938 -70076
rect 73014 -71258 73024 -70076
rect 72576 -71267 72658 -71262
rect 72932 -71263 73014 -71258
rect 73282 -71260 73292 -70078
rect 73368 -71260 73378 -70078
rect 73292 -71263 73374 -71260
rect 73632 -71262 73642 -70080
rect 73718 -71262 73728 -70080
rect 73994 -71262 74004 -70080
rect 74080 -71262 74090 -70080
rect 74346 -71256 74356 -70074
rect 74432 -71256 74442 -70074
rect 74356 -71261 74438 -71256
rect 73642 -71267 73724 -71262
rect 73998 -71263 74080 -71262
rect 74710 -71266 74720 -70084
rect 74796 -71266 74806 -70084
rect 75060 -71260 75070 -70078
rect 75146 -71260 75156 -70078
rect 75418 -71260 75428 -70078
rect 75504 -71260 75514 -70078
rect 75772 -71260 75782 -70078
rect 75858 -71260 75868 -70078
rect 76126 -71260 76136 -70078
rect 76212 -71260 76222 -70078
rect 76482 -71258 76492 -70076
rect 76568 -71258 76578 -70076
rect 75064 -71263 75146 -71260
rect 75422 -71261 75504 -71260
rect 75778 -71261 75860 -71260
rect 76136 -71263 76218 -71260
rect 76486 -71261 76568 -71258
rect 76844 -71270 76854 -70088
rect 76930 -71270 76940 -70088
rect 77188 -71262 77198 -70080
rect 77274 -71262 77284 -70080
rect 77544 -71262 77554 -70080
rect 77630 -71262 77640 -70080
rect 77908 -71256 77918 -70074
rect 77994 -71256 78004 -70074
rect 77916 -71259 77998 -71256
rect 77202 -71267 77284 -71262
rect 78262 -71266 78272 -70084
rect 78348 -71266 78358 -70084
rect 78624 -71262 78634 -70080
rect 78710 -71262 78720 -70080
rect 78982 -71262 78992 -70080
rect 79068 -71262 79078 -70080
rect 78986 -71263 79068 -71262
rect 79336 -71266 79346 -70084
rect 79422 -71266 79432 -70084
rect 79686 -71260 79696 -70078
rect 79772 -71260 79782 -70078
rect 79694 -71262 79704 -71260
rect 79766 -71262 79776 -71260
rect 79336 -71267 79418 -71266
rect 79694 -71267 79776 -71262
rect 80042 -71266 80052 -70084
rect 80128 -71266 80138 -70084
rect 80402 -71262 80412 -70080
rect 80488 -71262 80498 -70080
rect 80750 -71262 80760 -70080
rect 80836 -71262 80846 -70080
rect 81104 -71260 81114 -70078
rect 81190 -71260 81200 -70078
rect 81116 -71262 81126 -71260
rect 81188 -71262 81198 -71260
rect 80402 -71267 80484 -71262
rect 80758 -71263 80840 -71262
rect 81116 -71267 81198 -71262
rect 81468 -71266 81478 -70084
rect 81554 -71266 81564 -70084
rect 81820 -71262 81830 -70080
rect 81906 -71262 81916 -70080
rect 82166 -71262 82176 -70080
rect 82252 -71262 82262 -70080
rect 81826 -71267 81908 -71262
rect 82180 -71263 82262 -71262
rect 82524 -71268 82534 -70086
rect 82610 -71268 82620 -70086
rect 82884 -71266 82894 -70084
rect 82970 -71266 82980 -70084
rect 83254 -71256 83264 -70070
rect 83340 -71252 83350 -70070
rect 83326 -71256 83336 -71252
rect 83254 -71261 83336 -71256
rect 83606 -71268 83616 -70086
rect 83692 -71268 83702 -70086
rect 83970 -70113 83980 -70086
rect 83966 -70118 83980 -70113
rect 83966 -71262 83976 -70118
rect 83966 -71267 83980 -71262
rect 83970 -71268 83980 -71267
rect 84056 -71268 84066 -70086
rect 62348 -72616 62424 -71299
rect 62348 -72630 62426 -72616
rect 62710 -72630 62786 -71297
rect 63070 -72630 63146 -71285
rect 63414 -72630 63490 -71285
rect 63780 -72630 63856 -71283
rect 64134 -72630 64210 -71279
rect 56230 -73064 65354 -72630
rect 68302 -72676 68312 -71542
rect 68304 -72706 68314 -72676
rect 68376 -72706 68386 -71542
rect 68652 -72660 68662 -71526
rect 68654 -72684 68664 -72660
rect 68726 -72684 68736 -71526
rect 69008 -72660 69018 -71526
rect 69082 -72660 69092 -71526
rect 69366 -72660 69376 -71526
rect 68654 -72689 68736 -72684
rect 69368 -72684 69378 -72660
rect 69440 -72684 69450 -71526
rect 69714 -72664 69724 -71530
rect 69788 -72664 69798 -71530
rect 70078 -71531 70088 -71518
rect 70076 -71536 70088 -71531
rect 70076 -72646 70086 -71536
rect 70076 -72651 70088 -72646
rect 70078 -72652 70088 -72651
rect 70152 -72652 70162 -71518
rect 70440 -72660 70450 -71526
rect 70514 -72660 70524 -71526
rect 70780 -72664 70790 -71530
rect 70854 -72664 70864 -71530
rect 71138 -72672 71148 -71538
rect 71212 -72672 71222 -71538
rect 71494 -72664 71504 -71530
rect 71568 -72664 71578 -71530
rect 71848 -72660 71858 -71526
rect 71922 -72660 71932 -71526
rect 72208 -71541 72218 -71530
rect 72206 -71546 72218 -71541
rect 72206 -72656 72216 -71546
rect 72206 -72661 72218 -72656
rect 72208 -72664 72218 -72661
rect 72282 -72664 72292 -71530
rect 72562 -71539 72572 -71530
rect 72560 -71544 72572 -71539
rect 72560 -72654 72570 -71544
rect 72560 -72659 72572 -72654
rect 72562 -72664 72572 -72659
rect 72636 -72664 72646 -71530
rect 72934 -72664 72944 -71530
rect 73008 -72664 73018 -71530
rect 73276 -72676 73286 -71542
rect 73350 -72676 73360 -71542
rect 73632 -72660 73642 -71526
rect 73706 -72660 73716 -71526
rect 73978 -72652 73988 -71518
rect 74052 -72652 74062 -71518
rect 73978 -72657 74060 -72652
rect 73632 -72665 73714 -72660
rect 74342 -72672 74352 -71538
rect 74416 -72672 74426 -71538
rect 74704 -72666 74714 -71530
rect 74778 -72664 74788 -71530
rect 75060 -71567 75070 -71550
rect 75058 -71572 75070 -71567
rect 74776 -72666 74786 -72664
rect 74704 -72671 74786 -72666
rect 74342 -72675 74424 -72672
rect 69368 -72689 69450 -72684
rect 75058 -72682 75068 -71572
rect 75058 -72684 75070 -72682
rect 75134 -72684 75144 -71550
rect 75416 -72672 75426 -71538
rect 75490 -72672 75500 -71538
rect 75754 -72654 75764 -71518
rect 75828 -72652 75838 -71518
rect 76118 -72652 76128 -71518
rect 76192 -72652 76202 -71518
rect 75826 -72654 75836 -72652
rect 75754 -72659 75836 -72654
rect 76120 -72657 76202 -72652
rect 76468 -72652 76478 -71518
rect 76542 -72652 76552 -71518
rect 76468 -72657 76550 -72652
rect 76844 -72660 76854 -71526
rect 76918 -72660 76928 -71526
rect 77186 -72660 77196 -71526
rect 77260 -72660 77270 -71526
rect 77900 -71533 77910 -71514
rect 77898 -71538 77910 -71533
rect 76844 -72661 76926 -72660
rect 77186 -72665 77268 -72660
rect 77538 -72672 77548 -71538
rect 77612 -72672 77622 -71538
rect 77898 -72648 77908 -71538
rect 77974 -72648 77984 -71514
rect 77898 -72653 77980 -72648
rect 78264 -72652 78274 -71518
rect 78338 -72652 78348 -71518
rect 78264 -72655 78346 -72652
rect 78614 -72672 78624 -71538
rect 78688 -72672 78698 -71538
rect 75416 -72675 75498 -72672
rect 77538 -72677 77620 -72672
rect 78614 -72677 78696 -72672
rect 78978 -72676 78988 -71542
rect 79052 -72676 79062 -71542
rect 79328 -72652 79338 -71518
rect 79402 -72652 79412 -71518
rect 79684 -71545 79694 -71526
rect 79682 -71550 79694 -71545
rect 79328 -72657 79410 -72652
rect 79682 -72660 79692 -71550
rect 79758 -72660 79768 -71526
rect 79682 -72665 79764 -72660
rect 80036 -72664 80046 -71530
rect 80038 -72666 80048 -72664
rect 80110 -72666 80120 -71530
rect 80390 -71555 80400 -71538
rect 80038 -72671 80120 -72666
rect 80388 -71560 80400 -71555
rect 80388 -72670 80398 -71560
rect 80388 -72672 80400 -72670
rect 80464 -72672 80474 -71538
rect 80750 -72662 80760 -71526
rect 80824 -72660 80834 -71526
rect 81112 -71557 81122 -71538
rect 81110 -71562 81122 -71557
rect 80822 -72662 80832 -72660
rect 80750 -72667 80832 -72662
rect 81110 -72672 81120 -71562
rect 81186 -72672 81196 -71538
rect 81468 -72664 81478 -71530
rect 81542 -72664 81552 -71530
rect 81838 -72664 81848 -71530
rect 81912 -72664 81922 -71530
rect 81468 -72665 81550 -72664
rect 81838 -72667 81920 -72664
rect 82174 -72672 82184 -71538
rect 82248 -72672 82258 -71538
rect 80388 -72675 80470 -72672
rect 78980 -72677 79062 -72676
rect 81110 -72677 81192 -72672
rect 82176 -72675 82258 -72672
rect 82532 -72676 82542 -71542
rect 82606 -72676 82616 -71542
rect 82532 -72681 82614 -72676
rect 82896 -72684 82906 -71550
rect 82970 -71569 82980 -71550
rect 82970 -71574 82982 -71569
rect 82972 -72684 82982 -71574
rect 83246 -72664 83256 -71530
rect 83320 -72664 83330 -71530
rect 83248 -72667 83330 -72664
rect 75058 -72687 75140 -72684
rect 82900 -72689 82982 -72684
rect 83602 -72684 83612 -71550
rect 83676 -72684 83686 -71550
rect 83952 -72664 83962 -71530
rect 84026 -72664 84036 -71530
rect 83952 -72665 84034 -72664
rect 83602 -72689 83684 -72684
rect 68304 -72711 68386 -72706
rect 56842 -73396 56918 -73391
rect 56478 -73402 56554 -73397
rect 56842 -73402 56852 -73396
rect 56456 -73428 56488 -73402
rect 56544 -73428 56852 -73402
rect 56908 -73402 56918 -73396
rect 57546 -73402 57622 -73397
rect 58618 -73400 58694 -73395
rect 58618 -73402 58628 -73400
rect 56908 -73408 57556 -73402
rect 56908 -73428 57196 -73408
rect 57252 -73412 57556 -73408
rect 57612 -73408 58628 -73402
rect 57612 -73412 57916 -73408
rect 57252 -73428 57542 -73412
rect 56456 -74542 56466 -73428
rect 56560 -74534 56852 -73428
rect 56560 -74542 56854 -74534
rect 56948 -74542 57186 -73428
rect 57280 -74526 57542 -73428
rect 57636 -73422 57916 -73412
rect 57972 -73410 58628 -73408
rect 57972 -73412 58274 -73410
rect 58330 -73412 58628 -73410
rect 58684 -73402 58694 -73400
rect 58970 -73402 59046 -73399
rect 59332 -73400 59408 -73395
rect 59332 -73402 59342 -73400
rect 58684 -73404 59342 -73402
rect 58684 -73412 58980 -73404
rect 57972 -73422 58256 -73412
rect 57636 -74526 57890 -73422
rect 57280 -74540 57556 -74526
rect 57612 -74536 57890 -74526
rect 57984 -74526 58256 -73422
rect 58350 -74526 58616 -73412
rect 58710 -73428 58980 -73412
rect 59036 -73428 59342 -73404
rect 59398 -73402 59408 -73400
rect 59684 -73402 59760 -73399
rect 60754 -73402 60830 -73401
rect 61466 -73402 61542 -73399
rect 59398 -73404 64386 -73402
rect 59398 -73422 59694 -73404
rect 59750 -73406 61476 -73404
rect 59750 -73410 60764 -73406
rect 59750 -73412 60402 -73410
rect 59750 -73422 60052 -73412
rect 59398 -73428 59672 -73422
rect 58710 -74526 58970 -73428
rect 57984 -74536 58274 -74526
rect 57612 -74540 57916 -74536
rect 57280 -74542 57916 -74540
rect 56456 -74545 57196 -74542
rect 57186 -74546 57196 -74545
rect 57252 -74545 57916 -74542
rect 57252 -74546 57262 -74545
rect 57186 -74551 57262 -74546
rect 57906 -74546 57916 -74545
rect 57972 -74545 58274 -74536
rect 57972 -74546 57982 -74545
rect 57906 -74551 57982 -74546
rect 58264 -74548 58274 -74545
rect 58330 -74538 58628 -74526
rect 58684 -74538 58970 -74526
rect 58330 -74542 58970 -74538
rect 59064 -74542 59330 -73428
rect 59424 -74536 59672 -73428
rect 59766 -74536 60052 -73422
rect 59424 -74542 59694 -74536
rect 59750 -74542 60052 -74536
rect 58330 -74545 60052 -74542
rect 58330 -74548 58340 -74545
rect 58970 -74547 59046 -74545
rect 59684 -74547 59760 -74545
rect 58264 -74553 58340 -74548
rect 60042 -74550 60052 -74545
rect 60108 -74545 60402 -73412
rect 60108 -74550 60118 -74545
rect 60042 -74555 60118 -74550
rect 60392 -74548 60402 -74545
rect 60458 -74544 60764 -73410
rect 60820 -73410 61476 -73406
rect 60820 -74544 61118 -73410
rect 60458 -74545 61118 -74544
rect 60458 -74548 60468 -74545
rect 60392 -74553 60468 -74548
rect 60754 -74549 60830 -74545
rect 61108 -74548 61118 -74545
rect 61174 -74542 61476 -73410
rect 61532 -73408 64386 -73404
rect 61532 -73410 63966 -73408
rect 61532 -74542 61826 -73410
rect 61174 -74545 61826 -74542
rect 61174 -74548 61184 -74545
rect 61466 -74547 61542 -74545
rect 61108 -74553 61184 -74548
rect 61816 -74548 61826 -74545
rect 61882 -73414 62544 -73410
rect 61882 -74545 62188 -73414
rect 61882 -74548 61892 -74545
rect 61816 -74553 61892 -74548
rect 62178 -74552 62188 -74545
rect 62244 -74545 62544 -73414
rect 62244 -74552 62254 -74545
rect 62178 -74557 62254 -74552
rect 62534 -74548 62544 -74545
rect 62600 -73412 63966 -73410
rect 62600 -73414 63254 -73412
rect 62600 -74545 62894 -73414
rect 62600 -74548 62610 -74545
rect 62534 -74553 62610 -74548
rect 62884 -74552 62894 -74545
rect 62950 -74545 63254 -73414
rect 62950 -74552 62960 -74545
rect 62884 -74557 62960 -74552
rect 63244 -74550 63254 -74545
rect 63310 -73414 63966 -73412
rect 63310 -74545 63614 -73414
rect 63310 -74550 63320 -74545
rect 63244 -74555 63320 -74550
rect 63604 -74552 63614 -74545
rect 63670 -74545 63966 -73414
rect 63670 -74552 63680 -74545
rect 63956 -74546 63966 -74545
rect 64022 -74545 64320 -73408
rect 64022 -74546 64032 -74545
rect 63956 -74551 64032 -74546
rect 64310 -74546 64320 -74545
rect 64376 -74546 64386 -73408
rect 68052 -74360 84074 -73708
rect 64310 -74551 64386 -74546
rect 63604 -74557 63680 -74552
rect 56826 -74857 56902 -74853
rect 56458 -74858 64388 -74857
rect 56458 -74864 56836 -74858
rect 56458 -74874 56472 -74864
rect 56528 -74874 56836 -74864
rect 56892 -74862 64388 -74858
rect 56892 -74864 58612 -74862
rect 56892 -74870 57540 -74864
rect 56892 -74874 57180 -74870
rect 56458 -75988 56468 -74874
rect 56562 -75988 56828 -74874
rect 56922 -74884 57180 -74874
rect 57236 -74874 57540 -74870
rect 57596 -74868 58612 -74864
rect 58668 -74866 59326 -74862
rect 58668 -74868 58964 -74866
rect 57596 -74870 58600 -74868
rect 57596 -74874 57900 -74870
rect 57236 -74884 57532 -74874
rect 56922 -75988 57178 -74884
rect 56458 -76000 56472 -75988
rect 56462 -76002 56472 -76000
rect 56528 -75996 56836 -75988
rect 56892 -75996 57178 -75988
rect 56528 -75998 57178 -75996
rect 57272 -75988 57532 -74884
rect 57626 -74884 57900 -74874
rect 57956 -74872 58600 -74870
rect 57956 -74874 58258 -74872
rect 58314 -74874 58600 -74872
rect 57956 -74884 58246 -74874
rect 57626 -75988 57896 -74884
rect 57272 -75998 57540 -75988
rect 56528 -76000 57180 -75998
rect 56528 -76002 56538 -76000
rect 56826 -76001 56902 -76000
rect 56462 -76007 56538 -76002
rect 57170 -76008 57180 -76000
rect 57236 -76000 57540 -75998
rect 57236 -76008 57246 -76000
rect 57530 -76002 57540 -76000
rect 57596 -75998 57896 -75988
rect 57990 -75988 58246 -74884
rect 58340 -75982 58600 -74874
rect 58694 -74874 58964 -74868
rect 59020 -74868 59326 -74866
rect 59382 -74866 64388 -74862
rect 59382 -74868 59678 -74866
rect 59020 -74874 59320 -74868
rect 58694 -75982 58960 -74874
rect 58340 -75988 58612 -75982
rect 57990 -75998 58258 -75988
rect 57596 -76000 57900 -75998
rect 57596 -76002 57606 -76000
rect 57530 -76007 57606 -76002
rect 57170 -76013 57246 -76008
rect 57890 -76008 57900 -76000
rect 57956 -76000 58258 -75998
rect 57956 -76008 57966 -76000
rect 57890 -76013 57966 -76008
rect 58248 -76010 58258 -76000
rect 58314 -76000 58612 -75988
rect 58668 -75988 58960 -75982
rect 59054 -75982 59320 -74874
rect 59414 -74884 59678 -74868
rect 59734 -74868 61460 -74866
rect 59734 -74872 60748 -74868
rect 59734 -74874 60386 -74872
rect 59734 -74884 60036 -74874
rect 59414 -75982 59668 -74884
rect 59054 -75988 59326 -75982
rect 58668 -76000 58964 -75988
rect 58314 -76010 58324 -76000
rect 58602 -76005 58678 -76000
rect 58954 -76004 58964 -76000
rect 59020 -76000 59326 -75988
rect 59382 -75998 59668 -75982
rect 59762 -75998 60036 -74884
rect 59382 -76000 59678 -75998
rect 59020 -76004 59030 -76000
rect 58954 -76009 59030 -76004
rect 59316 -76005 59392 -76000
rect 59668 -76004 59678 -76000
rect 59734 -76000 60036 -75998
rect 59734 -76004 59744 -76000
rect 59668 -76009 59744 -76004
rect 58248 -76015 58324 -76010
rect 60026 -76012 60036 -76000
rect 60092 -76000 60386 -74874
rect 60092 -76012 60102 -76000
rect 60026 -76017 60102 -76012
rect 60376 -76010 60386 -76000
rect 60442 -76000 60748 -74872
rect 60442 -76010 60452 -76000
rect 60376 -76015 60452 -76010
rect 60738 -76006 60748 -76000
rect 60804 -74872 61460 -74868
rect 60804 -76000 61102 -74872
rect 60804 -76006 60814 -76000
rect 60738 -76011 60814 -76006
rect 61092 -76010 61102 -76000
rect 61158 -76000 61460 -74872
rect 61158 -76010 61168 -76000
rect 61450 -76004 61460 -76000
rect 61516 -74870 64388 -74866
rect 61516 -74872 63950 -74870
rect 61516 -76000 61810 -74872
rect 61516 -76004 61526 -76000
rect 61450 -76009 61526 -76004
rect 61092 -76015 61168 -76010
rect 61800 -76010 61810 -76000
rect 61866 -74876 62528 -74872
rect 61866 -76000 62172 -74876
rect 61866 -76010 61876 -76000
rect 61800 -76015 61876 -76010
rect 62162 -76014 62172 -76000
rect 62228 -76000 62528 -74876
rect 62228 -76014 62238 -76000
rect 62162 -76019 62238 -76014
rect 62518 -76010 62528 -76000
rect 62584 -74874 63950 -74872
rect 62584 -74876 63238 -74874
rect 62584 -76000 62878 -74876
rect 62584 -76010 62594 -76000
rect 62518 -76015 62594 -76010
rect 62868 -76014 62878 -76000
rect 62934 -76000 63238 -74876
rect 62934 -76014 62944 -76000
rect 62868 -76019 62944 -76014
rect 63228 -76012 63238 -76000
rect 63294 -74876 63950 -74874
rect 63294 -76000 63598 -74876
rect 63294 -76012 63304 -76000
rect 63228 -76017 63304 -76012
rect 63588 -76014 63598 -76000
rect 63654 -76000 63950 -74876
rect 63654 -76014 63664 -76000
rect 63940 -76008 63950 -76000
rect 64006 -76000 64304 -74870
rect 64006 -76008 64016 -76000
rect 63940 -76013 64016 -76008
rect 64294 -76008 64304 -76000
rect 64360 -76000 64388 -74870
rect 64360 -76008 64370 -76000
rect 64294 -76013 64370 -76008
rect 63588 -76019 63664 -76014
rect 56832 -77246 56908 -77241
rect 56468 -77252 56544 -77247
rect 56468 -77255 56478 -77252
rect 56446 -77284 56478 -77255
rect 56534 -77255 56544 -77252
rect 56832 -77255 56842 -77246
rect 56534 -77284 56842 -77255
rect 56898 -77255 56908 -77246
rect 57536 -77252 57612 -77247
rect 57176 -77255 57252 -77253
rect 57536 -77255 57546 -77252
rect 56898 -77258 57546 -77255
rect 56898 -77284 57186 -77258
rect 56446 -78398 56456 -77284
rect 56550 -78398 56816 -77284
rect 56910 -77294 57186 -77284
rect 57242 -77284 57546 -77258
rect 57602 -77255 57612 -77252
rect 58608 -77250 58684 -77245
rect 57896 -77255 57972 -77253
rect 58608 -77255 58618 -77250
rect 57602 -77258 58618 -77255
rect 57602 -77284 57906 -77258
rect 57242 -77294 57520 -77284
rect 56910 -78398 57166 -77294
rect 57156 -78408 57166 -78398
rect 57260 -78398 57520 -77294
rect 57614 -77294 57906 -77284
rect 57962 -77260 58618 -77258
rect 57962 -77284 58264 -77260
rect 58320 -77278 58618 -77260
rect 58674 -77255 58684 -77250
rect 58960 -77254 59036 -77249
rect 58960 -77255 58970 -77254
rect 58674 -77278 58970 -77255
rect 58320 -77284 58588 -77278
rect 57962 -77294 58234 -77284
rect 57614 -78398 57884 -77294
rect 57260 -78408 57270 -78398
rect 57874 -78408 57884 -78398
rect 57978 -78398 58234 -77294
rect 58328 -78392 58588 -77284
rect 58682 -77284 58970 -77278
rect 59026 -77255 59036 -77254
rect 59322 -77250 59398 -77245
rect 59322 -77255 59332 -77250
rect 59026 -77278 59332 -77255
rect 59388 -77255 59398 -77250
rect 59674 -77254 59750 -77249
rect 59674 -77255 59684 -77254
rect 59388 -77278 59684 -77255
rect 59026 -77284 59308 -77278
rect 58682 -78392 58948 -77284
rect 59042 -78392 59308 -77284
rect 59402 -77294 59684 -77278
rect 59740 -77255 59750 -77254
rect 60744 -77255 60820 -77251
rect 61456 -77254 61532 -77249
rect 61456 -77255 61466 -77254
rect 59740 -77256 61466 -77255
rect 59740 -77260 60754 -77256
rect 59740 -77262 60392 -77260
rect 59740 -77294 60042 -77262
rect 59402 -78392 59656 -77294
rect 58328 -78398 58948 -78392
rect 59042 -78398 59656 -78392
rect 57978 -78408 57988 -78398
rect 58254 -78403 58330 -78398
rect 59646 -78408 59656 -78398
rect 59750 -78398 60042 -77294
rect 59750 -78408 59760 -78398
rect 60032 -78400 60042 -78398
rect 60098 -78398 60392 -77262
rect 60448 -78394 60754 -77260
rect 60810 -77260 61466 -77256
rect 60810 -78394 61108 -77260
rect 60448 -78398 61108 -78394
rect 61164 -78392 61466 -77260
rect 61522 -77255 61532 -77254
rect 63946 -77255 64022 -77253
rect 64300 -77255 64376 -77253
rect 61522 -77258 64376 -77255
rect 61522 -77260 63956 -77258
rect 61522 -78392 61816 -77260
rect 61164 -78398 61816 -78392
rect 61872 -77264 62534 -77260
rect 61872 -78398 62178 -77264
rect 60098 -78400 60108 -78398
rect 60032 -78405 60108 -78400
rect 60382 -78403 60458 -78398
rect 60744 -78399 60820 -78398
rect 61098 -78403 61174 -78398
rect 61806 -78403 61882 -78398
rect 62168 -78402 62178 -78398
rect 62234 -78398 62534 -77264
rect 62590 -77262 63956 -77260
rect 62590 -77264 63244 -77262
rect 62590 -78398 62884 -77264
rect 62234 -78402 62244 -78398
rect 62168 -78407 62244 -78402
rect 62524 -78403 62600 -78398
rect 62874 -78402 62884 -78398
rect 62940 -78398 63244 -77264
rect 62940 -78402 62950 -78398
rect 62874 -78407 62950 -78402
rect 63234 -78400 63244 -78398
rect 63300 -77264 63956 -77262
rect 63300 -78398 63604 -77264
rect 63300 -78400 63310 -78398
rect 63234 -78405 63310 -78400
rect 63594 -78402 63604 -78398
rect 63660 -78396 63956 -77264
rect 64012 -78396 64310 -77258
rect 64366 -78396 64376 -77258
rect 63660 -78398 64376 -78396
rect 63660 -78402 63670 -78398
rect 63946 -78401 64022 -78398
rect 64300 -78401 64376 -78398
rect 63594 -78407 63670 -78402
rect 56816 -78708 56892 -78703
rect 56816 -78709 56826 -78708
rect 56430 -78714 56826 -78709
rect 56430 -78720 56462 -78714
rect 56518 -78720 56826 -78714
rect 56882 -78709 56892 -78708
rect 58592 -78709 58668 -78707
rect 59306 -78709 59382 -78707
rect 56882 -78712 64360 -78709
rect 56882 -78714 58602 -78712
rect 58658 -78714 59316 -78712
rect 59372 -78714 64360 -78712
rect 56882 -78720 57530 -78714
rect 57586 -78720 58572 -78714
rect 56430 -79834 56440 -78720
rect 56534 -79834 56800 -78720
rect 56894 -78730 57170 -78720
rect 57226 -78730 57504 -78720
rect 56894 -79834 57150 -78730
rect 56430 -79852 56462 -79834
rect 56518 -79846 56826 -79834
rect 56882 -79844 57150 -79834
rect 57244 -79834 57504 -78730
rect 57598 -78730 57890 -78720
rect 57946 -78730 58218 -78720
rect 57598 -79834 57868 -78730
rect 57244 -79844 57530 -79834
rect 56882 -79846 57170 -79844
rect 56518 -79852 57170 -79846
rect 56452 -79857 56528 -79852
rect 57160 -79858 57170 -79852
rect 57226 -79852 57530 -79844
rect 57586 -79844 57868 -79834
rect 57962 -79834 58218 -78730
rect 58312 -79828 58572 -78720
rect 58666 -78716 59292 -78714
rect 58666 -78720 58954 -78716
rect 59010 -78720 59292 -78716
rect 58666 -79828 58932 -78720
rect 58312 -79834 58602 -79828
rect 57962 -79844 58248 -79834
rect 57586 -79852 57890 -79844
rect 57226 -79858 57236 -79852
rect 57520 -79857 57596 -79852
rect 57160 -79863 57236 -79858
rect 57880 -79858 57890 -79852
rect 57946 -79852 58248 -79844
rect 57946 -79858 57956 -79852
rect 57880 -79863 57956 -79858
rect 58238 -79860 58248 -79852
rect 58304 -79850 58602 -79834
rect 58658 -79834 58932 -79828
rect 59026 -79828 59292 -78720
rect 59386 -78716 64360 -78714
rect 59386 -78730 59668 -78716
rect 59724 -78718 61450 -78716
rect 59724 -78722 60738 -78718
rect 59724 -78724 60376 -78722
rect 59724 -78730 60026 -78724
rect 59386 -79828 59640 -78730
rect 59026 -79834 59316 -79828
rect 58658 -79850 58954 -79834
rect 58304 -79852 58954 -79850
rect 58304 -79860 58314 -79852
rect 58592 -79855 58668 -79852
rect 58944 -79854 58954 -79852
rect 59010 -79850 59316 -79834
rect 59372 -79844 59640 -79828
rect 59734 -79844 60026 -78730
rect 59372 -79850 59668 -79844
rect 59010 -79852 59668 -79850
rect 59010 -79854 59020 -79852
rect 58944 -79859 59020 -79854
rect 59306 -79855 59382 -79852
rect 59658 -79854 59668 -79852
rect 59724 -79852 60026 -79844
rect 59724 -79854 59734 -79852
rect 59658 -79859 59734 -79854
rect 58238 -79865 58314 -79860
rect 60016 -79862 60026 -79852
rect 60082 -79852 60376 -78724
rect 60082 -79862 60092 -79852
rect 60016 -79867 60092 -79862
rect 60366 -79860 60376 -79852
rect 60432 -79852 60738 -78722
rect 60432 -79860 60442 -79852
rect 60366 -79865 60442 -79860
rect 60728 -79856 60738 -79852
rect 60794 -78722 61450 -78718
rect 60794 -79852 61092 -78722
rect 60794 -79856 60804 -79852
rect 60728 -79861 60804 -79856
rect 61082 -79860 61092 -79852
rect 61148 -79852 61450 -78722
rect 61148 -79860 61158 -79852
rect 61440 -79854 61450 -79852
rect 61506 -78720 64360 -78716
rect 61506 -78722 63940 -78720
rect 61506 -79852 61800 -78722
rect 61506 -79854 61516 -79852
rect 61440 -79859 61516 -79854
rect 61082 -79865 61158 -79860
rect 61790 -79860 61800 -79852
rect 61856 -78726 62518 -78722
rect 61856 -79852 62162 -78726
rect 61856 -79860 61866 -79852
rect 61790 -79865 61866 -79860
rect 62152 -79864 62162 -79852
rect 62218 -79852 62518 -78726
rect 62218 -79864 62228 -79852
rect 62152 -79869 62228 -79864
rect 62508 -79860 62518 -79852
rect 62574 -78724 63940 -78722
rect 62574 -78726 63228 -78724
rect 62574 -79852 62868 -78726
rect 62574 -79860 62584 -79852
rect 62508 -79865 62584 -79860
rect 62858 -79864 62868 -79852
rect 62924 -79852 63228 -78726
rect 62924 -79864 62934 -79852
rect 62858 -79869 62934 -79864
rect 63218 -79862 63228 -79852
rect 63284 -78726 63940 -78724
rect 63284 -79852 63588 -78726
rect 63284 -79862 63294 -79852
rect 63218 -79867 63294 -79862
rect 63578 -79864 63588 -79852
rect 63644 -79852 63940 -78726
rect 63644 -79864 63654 -79852
rect 63930 -79858 63940 -79852
rect 63996 -79852 64294 -78720
rect 63996 -79858 64006 -79852
rect 63930 -79863 64006 -79858
rect 64284 -79858 64294 -79852
rect 64350 -79858 64360 -78720
rect 64284 -79863 64360 -79858
rect 63578 -79869 63654 -79864
rect 67376 -80074 80234 -79244
rect 56842 -81212 56918 -81207
rect 56478 -81218 56554 -81213
rect 56842 -81218 56852 -81212
rect 56478 -82356 56488 -81218
rect 56544 -82350 56852 -81218
rect 56908 -81218 56918 -81212
rect 57546 -81218 57622 -81213
rect 58618 -81216 58694 -81211
rect 58618 -81218 58628 -81216
rect 56908 -81224 57556 -81218
rect 56908 -82350 57196 -81224
rect 56544 -82356 57196 -82350
rect 56478 -82361 57196 -82356
rect 57186 -82362 57196 -82361
rect 57252 -82356 57556 -81224
rect 57612 -81224 58628 -81218
rect 57612 -82356 57916 -81224
rect 57252 -82361 57916 -82356
rect 57252 -82362 57262 -82361
rect 57186 -82367 57262 -82362
rect 57906 -82362 57916 -82361
rect 57972 -81226 58628 -81224
rect 57972 -82361 58274 -81226
rect 57972 -82362 57982 -82361
rect 57906 -82367 57982 -82362
rect 58264 -82364 58274 -82361
rect 58330 -82354 58628 -81226
rect 58684 -81218 58694 -81216
rect 58970 -81218 59046 -81215
rect 59332 -81216 59408 -81211
rect 59332 -81218 59342 -81216
rect 58684 -81220 59342 -81218
rect 58684 -82354 58980 -81220
rect 58330 -82358 58980 -82354
rect 59036 -82354 59342 -81220
rect 59398 -81218 59408 -81216
rect 59684 -81218 59760 -81215
rect 60754 -81218 60830 -81217
rect 61466 -81218 61542 -81215
rect 59398 -81220 64408 -81218
rect 59398 -82354 59694 -81220
rect 59036 -82358 59694 -82354
rect 59750 -81222 61476 -81220
rect 59750 -81226 60764 -81222
rect 59750 -81228 60402 -81226
rect 59750 -82358 60052 -81228
rect 58330 -82361 60052 -82358
rect 58330 -82364 58340 -82361
rect 58970 -82363 59046 -82361
rect 59684 -82363 59760 -82361
rect 58264 -82369 58340 -82364
rect 60042 -82366 60052 -82361
rect 60108 -82361 60402 -81228
rect 60108 -82366 60118 -82361
rect 60042 -82371 60118 -82366
rect 60392 -82364 60402 -82361
rect 60458 -82360 60764 -81226
rect 60820 -81226 61476 -81222
rect 60820 -81246 61118 -81226
rect 61174 -81230 61476 -81226
rect 61532 -81224 64408 -81220
rect 61532 -81226 63966 -81224
rect 61532 -81230 61826 -81226
rect 61882 -81230 62544 -81226
rect 61174 -81246 61462 -81230
rect 60820 -82360 61102 -81246
rect 61196 -82344 61462 -81246
rect 61556 -82344 61810 -81230
rect 61904 -82344 62170 -81230
rect 62264 -81236 62544 -81230
rect 62600 -81228 63966 -81226
rect 62600 -81230 63254 -81228
rect 62600 -81236 62894 -81230
rect 62950 -81236 63254 -81230
rect 63310 -81230 63966 -81228
rect 64022 -81230 64320 -81224
rect 64376 -81230 64408 -81224
rect 63310 -81236 63614 -81230
rect 62264 -82344 62530 -81236
rect 61196 -82358 61476 -82344
rect 61532 -82358 61826 -82344
rect 61196 -82360 61826 -82358
rect 60458 -82361 61118 -82360
rect 60458 -82364 60468 -82361
rect 60392 -82369 60468 -82364
rect 60754 -82365 60830 -82361
rect 61108 -82364 61118 -82361
rect 61174 -82361 61826 -82360
rect 61174 -82364 61184 -82361
rect 61466 -82363 61542 -82361
rect 61108 -82369 61184 -82364
rect 61816 -82364 61826 -82361
rect 61882 -82361 62188 -82344
rect 61882 -82364 61892 -82361
rect 61816 -82369 61892 -82364
rect 62178 -82368 62188 -82361
rect 62244 -82350 62530 -82344
rect 62624 -82350 62884 -81236
rect 62978 -82350 63234 -81236
rect 63328 -81246 63614 -81236
rect 63670 -81246 63952 -81230
rect 63328 -82350 63594 -81246
rect 62244 -82361 62544 -82350
rect 62244 -82368 62254 -82361
rect 62178 -82373 62254 -82368
rect 62534 -82364 62544 -82361
rect 62600 -82361 62894 -82350
rect 62600 -82364 62610 -82361
rect 62534 -82369 62610 -82364
rect 62884 -82368 62894 -82361
rect 62950 -82361 63254 -82350
rect 62950 -82368 62960 -82361
rect 62884 -82373 62960 -82368
rect 63244 -82366 63254 -82361
rect 63310 -82360 63594 -82350
rect 63688 -82344 63952 -81246
rect 64046 -82344 64296 -81230
rect 64390 -82344 64408 -81230
rect 63688 -82360 63966 -82344
rect 63310 -82361 63614 -82360
rect 63310 -82366 63320 -82361
rect 63244 -82371 63320 -82366
rect 63604 -82368 63614 -82361
rect 63670 -82361 63966 -82360
rect 63670 -82368 63680 -82361
rect 63956 -82362 63966 -82361
rect 64022 -82361 64320 -82344
rect 64022 -82362 64032 -82361
rect 63956 -82367 64032 -82362
rect 64310 -82362 64320 -82361
rect 64376 -82361 64408 -82344
rect 64376 -82362 64386 -82361
rect 64310 -82367 64386 -82362
rect 63604 -82373 63680 -82368
rect 56826 -82674 56902 -82669
rect 56462 -82680 56538 -82675
rect 56462 -83818 56472 -82680
rect 56528 -82681 56538 -82680
rect 56826 -82681 56836 -82674
rect 56528 -83812 56836 -82681
rect 56892 -82681 56902 -82674
rect 57530 -82680 57606 -82675
rect 57530 -82681 57540 -82680
rect 56892 -82686 57540 -82681
rect 56892 -83812 57180 -82686
rect 56528 -83818 57180 -83812
rect 56462 -83823 57180 -83818
rect 56463 -83824 57180 -83823
rect 57236 -83818 57540 -82686
rect 57596 -82681 57606 -82680
rect 58602 -82678 58678 -82673
rect 58602 -82681 58612 -82678
rect 57596 -82686 58612 -82681
rect 57596 -83818 57900 -82686
rect 57236 -83824 57900 -83818
rect 57956 -82688 58612 -82686
rect 57956 -83824 58258 -82688
rect 57170 -83829 57246 -83824
rect 57890 -83829 57966 -83824
rect 58248 -83826 58258 -83824
rect 58314 -83816 58612 -82688
rect 58668 -82681 58678 -82678
rect 58954 -82681 59030 -82677
rect 59316 -82678 59392 -82673
rect 59316 -82681 59326 -82678
rect 58668 -82682 59326 -82681
rect 58668 -83816 58964 -82682
rect 58314 -83820 58964 -83816
rect 59020 -83816 59326 -82682
rect 59382 -82681 59392 -82678
rect 59668 -82681 59744 -82677
rect 60738 -82681 60814 -82679
rect 61434 -82681 61444 -82676
rect 59382 -82682 61444 -82681
rect 61538 -82681 61548 -82676
rect 61778 -82681 61788 -82676
rect 59382 -83816 59678 -82682
rect 59020 -83820 59678 -83816
rect 59734 -82684 61444 -82682
rect 59734 -82688 60748 -82684
rect 59734 -82690 60386 -82688
rect 59734 -83820 60036 -82690
rect 58314 -83824 60036 -83820
rect 58314 -83826 58324 -83824
rect 58954 -83825 59030 -83824
rect 59668 -83825 59744 -83824
rect 58248 -83831 58324 -83826
rect 60026 -83828 60036 -83824
rect 60092 -83824 60386 -82690
rect 60092 -83828 60102 -83824
rect 60026 -83833 60102 -83828
rect 60376 -83826 60386 -83824
rect 60442 -83822 60748 -82688
rect 60804 -82688 61444 -82684
rect 60804 -82702 61102 -82688
rect 61158 -82702 61444 -82688
rect 60804 -83816 61086 -82702
rect 61180 -83790 61444 -82702
rect 61538 -83790 61788 -82681
rect 61882 -82681 61892 -82676
rect 62154 -82681 62164 -82676
rect 61882 -83790 62164 -82681
rect 62258 -82681 62268 -82676
rect 62504 -82681 62514 -82676
rect 62258 -83790 62514 -82681
rect 62608 -82681 62618 -82676
rect 63566 -82681 63576 -82670
rect 62608 -82686 63576 -82681
rect 62608 -83790 62856 -82686
rect 62950 -82690 63576 -82686
rect 62950 -82692 63238 -82690
rect 63294 -82692 63576 -82690
rect 63670 -82681 63680 -82670
rect 63670 -82686 64393 -82681
rect 61180 -83816 61460 -83790
rect 60804 -83822 61102 -83816
rect 60442 -83824 61102 -83822
rect 60442 -83826 60452 -83824
rect 60376 -83831 60452 -83826
rect 60738 -83827 60814 -83824
rect 61092 -83826 61102 -83824
rect 61158 -83820 61460 -83816
rect 61516 -83820 61810 -83790
rect 61158 -83824 61810 -83820
rect 61158 -83826 61168 -83824
rect 61450 -83825 61526 -83824
rect 61092 -83831 61168 -83826
rect 61800 -83826 61810 -83824
rect 61866 -83824 62172 -83790
rect 61866 -83826 61876 -83824
rect 61800 -83831 61876 -83826
rect 62162 -83830 62172 -83824
rect 62228 -83824 62528 -83790
rect 62228 -83830 62238 -83824
rect 62162 -83835 62238 -83830
rect 62518 -83826 62528 -83824
rect 62584 -83800 62856 -83790
rect 62950 -83800 63216 -82692
rect 62584 -83824 62878 -83800
rect 62584 -83826 62594 -83824
rect 62518 -83831 62594 -83826
rect 62868 -83830 62878 -83824
rect 62934 -83806 63216 -83800
rect 63310 -83784 63576 -82692
rect 63670 -83784 63920 -82686
rect 63310 -83806 63598 -83784
rect 62934 -83824 63238 -83806
rect 62934 -83830 62944 -83824
rect 62868 -83835 62944 -83830
rect 63228 -83828 63238 -83824
rect 63294 -83824 63598 -83806
rect 63294 -83828 63304 -83824
rect 63228 -83833 63304 -83828
rect 63588 -83830 63598 -83824
rect 63654 -83800 63920 -83784
rect 64014 -82692 64304 -82686
rect 64360 -82692 64393 -82686
rect 64014 -83800 64286 -82692
rect 63654 -83824 63950 -83800
rect 64006 -83806 64286 -83800
rect 64380 -83806 64393 -82692
rect 64006 -83824 64304 -83806
rect 64360 -83824 64393 -83806
rect 63654 -83830 63664 -83824
rect 63940 -83829 64016 -83824
rect 64294 -83829 64370 -83824
rect 63588 -83835 63664 -83830
rect 56814 -85032 56890 -85027
rect 56450 -85038 56526 -85033
rect 56450 -86176 56460 -85038
rect 56516 -85039 56526 -85038
rect 56814 -85039 56824 -85032
rect 56516 -86170 56824 -85039
rect 56880 -85039 56890 -85032
rect 57518 -85038 57594 -85033
rect 57518 -85039 57528 -85038
rect 56880 -85044 57528 -85039
rect 56880 -86170 57168 -85044
rect 56516 -86176 57168 -86170
rect 56450 -86182 57168 -86176
rect 57224 -86176 57528 -85044
rect 57584 -85039 57594 -85038
rect 58590 -85036 58666 -85031
rect 58590 -85039 58600 -85036
rect 57584 -85044 58600 -85039
rect 57584 -86176 57888 -85044
rect 57224 -86182 57888 -86176
rect 57944 -85046 58600 -85044
rect 57944 -86182 58246 -85046
rect 57158 -86187 57234 -86182
rect 57878 -86187 57954 -86182
rect 58236 -86184 58246 -86182
rect 58302 -86174 58600 -85046
rect 58656 -85039 58666 -85036
rect 58942 -85039 59018 -85035
rect 59304 -85036 59380 -85031
rect 59304 -85039 59314 -85036
rect 58656 -85040 59314 -85039
rect 58656 -86174 58952 -85040
rect 58302 -86178 58952 -86174
rect 59008 -86174 59314 -85040
rect 59370 -85039 59380 -85036
rect 59656 -85039 59732 -85035
rect 60726 -85039 60802 -85037
rect 61438 -85039 61514 -85035
rect 61768 -85039 61778 -85036
rect 59370 -85040 61778 -85039
rect 59370 -86174 59666 -85040
rect 59008 -86178 59666 -86174
rect 59722 -85042 61448 -85040
rect 59722 -85046 60736 -85042
rect 59722 -85048 60374 -85046
rect 59722 -86178 60024 -85048
rect 58302 -86182 60024 -86178
rect 58302 -86184 58312 -86182
rect 58942 -86183 59018 -86182
rect 59656 -86183 59732 -86182
rect 58236 -86189 58312 -86184
rect 60014 -86186 60024 -86182
rect 60080 -86182 60374 -85048
rect 60080 -86186 60090 -86182
rect 60014 -86191 60090 -86186
rect 60364 -86184 60374 -86182
rect 60430 -86180 60736 -85046
rect 60792 -85046 61448 -85042
rect 61504 -85046 61778 -85040
rect 61872 -85039 61882 -85036
rect 62144 -85039 62154 -85036
rect 60792 -85068 61090 -85046
rect 61146 -85068 61418 -85046
rect 60792 -86180 61068 -85068
rect 60430 -86182 61068 -86180
rect 61162 -86160 61418 -85068
rect 61512 -86150 61778 -85046
rect 61872 -86150 62154 -85039
rect 62248 -85039 62258 -85036
rect 62482 -85039 62492 -85036
rect 62248 -86150 62492 -85039
rect 62586 -85039 62596 -85036
rect 64260 -85039 64270 -85024
rect 62586 -85044 64270 -85039
rect 64364 -85039 64374 -85024
rect 62586 -85048 63938 -85044
rect 62586 -85050 63226 -85048
rect 62586 -85064 62866 -85050
rect 62922 -85064 63226 -85050
rect 63282 -85050 63938 -85048
rect 63282 -85052 63586 -85050
rect 63642 -85052 63938 -85050
rect 63994 -85052 64270 -85044
rect 63282 -85064 63566 -85052
rect 62586 -86150 62840 -85064
rect 61512 -86160 61798 -86150
rect 61162 -86178 61448 -86160
rect 61504 -86178 61798 -86160
rect 61162 -86182 61798 -86178
rect 60430 -86184 60440 -86182
rect 60364 -86189 60440 -86184
rect 60726 -86185 60802 -86182
rect 61080 -86184 61090 -86182
rect 61146 -86184 61156 -86182
rect 61438 -86183 61514 -86182
rect 61080 -86189 61156 -86184
rect 61788 -86184 61798 -86182
rect 61854 -86182 62160 -86150
rect 61854 -86184 61864 -86182
rect 61788 -86189 61864 -86184
rect 62150 -86188 62160 -86182
rect 62216 -86182 62516 -86150
rect 62216 -86188 62226 -86182
rect 62150 -86193 62226 -86188
rect 62506 -86184 62516 -86182
rect 62572 -86178 62840 -86150
rect 62934 -86178 63206 -85064
rect 63300 -86166 63566 -85064
rect 63660 -86166 63926 -85052
rect 64020 -86138 64270 -85052
rect 64364 -86138 64380 -85039
rect 64020 -86166 64292 -86138
rect 63300 -86178 63586 -86166
rect 62572 -86182 62866 -86178
rect 62572 -86184 62582 -86182
rect 62506 -86189 62582 -86184
rect 62856 -86188 62866 -86182
rect 62922 -86182 63226 -86178
rect 62922 -86188 62932 -86182
rect 62856 -86193 62932 -86188
rect 63216 -86186 63226 -86182
rect 63282 -86182 63586 -86178
rect 63282 -86186 63292 -86182
rect 63216 -86191 63292 -86186
rect 63576 -86188 63586 -86182
rect 63642 -86182 63938 -86166
rect 63994 -86182 64292 -86166
rect 64348 -86182 64380 -86138
rect 63642 -86188 63652 -86182
rect 63928 -86187 64004 -86182
rect 64282 -86187 64358 -86182
rect 63576 -86193 63652 -86188
rect 56798 -86494 56874 -86489
rect 56434 -86500 56510 -86495
rect 56798 -86500 56808 -86494
rect 56434 -87638 56444 -86500
rect 56500 -87632 56808 -86500
rect 56864 -86500 56874 -86494
rect 57502 -86500 57578 -86495
rect 58574 -86498 58650 -86493
rect 58574 -86500 58584 -86498
rect 56864 -86506 57512 -86500
rect 56864 -87632 57152 -86506
rect 56500 -87638 57152 -87632
rect 56434 -87643 57152 -87638
rect 57142 -87644 57152 -87643
rect 57208 -87638 57512 -86506
rect 57568 -86506 58584 -86500
rect 57568 -87638 57872 -86506
rect 57208 -87643 57872 -87638
rect 57208 -87644 57218 -87643
rect 57142 -87649 57218 -87644
rect 57862 -87644 57872 -87643
rect 57928 -86508 58584 -86506
rect 57928 -87643 58230 -86508
rect 57928 -87644 57938 -87643
rect 57862 -87649 57938 -87644
rect 58220 -87646 58230 -87643
rect 58286 -87636 58584 -86508
rect 58640 -86500 58650 -86498
rect 58926 -86500 59002 -86497
rect 59288 -86498 59364 -86493
rect 59288 -86500 59298 -86498
rect 58640 -86502 59298 -86500
rect 58640 -87636 58936 -86502
rect 58286 -87640 58936 -87636
rect 58992 -87636 59298 -86502
rect 59354 -86500 59364 -86498
rect 59640 -86500 59716 -86497
rect 60710 -86500 60786 -86499
rect 61048 -86500 61058 -86480
rect 59354 -86502 61058 -86500
rect 59354 -87636 59650 -86502
rect 58992 -87640 59650 -87636
rect 59706 -86504 61058 -86502
rect 59706 -86508 60720 -86504
rect 59706 -86510 60358 -86508
rect 59706 -87640 60008 -86510
rect 58286 -87643 60008 -87640
rect 58286 -87646 58296 -87643
rect 58926 -87645 59002 -87643
rect 59640 -87645 59716 -87643
rect 58220 -87651 58296 -87646
rect 59998 -87648 60008 -87643
rect 60064 -87643 60358 -86510
rect 60064 -87648 60074 -87643
rect 59998 -87653 60074 -87648
rect 60348 -87646 60358 -87643
rect 60414 -87642 60720 -86508
rect 60776 -87594 61058 -86504
rect 61152 -86500 61162 -86480
rect 61422 -86498 61498 -86497
rect 61408 -86500 61418 -86498
rect 61152 -87594 61418 -86500
rect 61512 -86500 61522 -86498
rect 62122 -86500 62132 -86498
rect 60776 -87642 61074 -87594
rect 60414 -87643 61074 -87642
rect 60414 -87646 60424 -87643
rect 60348 -87651 60424 -87646
rect 60710 -87647 60786 -87643
rect 61064 -87646 61074 -87643
rect 61130 -87612 61418 -87594
rect 61512 -86508 62132 -86500
rect 61512 -86518 61782 -86508
rect 61838 -86518 62132 -86508
rect 62226 -86500 62236 -86498
rect 62482 -86500 62492 -86492
rect 61512 -87612 61772 -86518
rect 61130 -87640 61432 -87612
rect 61488 -87632 61772 -87612
rect 61866 -87612 62132 -86518
rect 62226 -87606 62492 -86500
rect 62586 -86500 62596 -86492
rect 63550 -86500 63560 -86498
rect 62586 -86508 63560 -86500
rect 62586 -86512 63200 -86508
rect 62586 -86518 62850 -86512
rect 62906 -86518 63200 -86512
rect 62586 -87606 62840 -86518
rect 62226 -87612 62500 -87606
rect 61866 -87632 62144 -87612
rect 61488 -87640 61782 -87632
rect 61130 -87643 61782 -87640
rect 61130 -87646 61140 -87643
rect 61422 -87645 61498 -87643
rect 61064 -87651 61140 -87646
rect 61772 -87646 61782 -87643
rect 61838 -87643 62144 -87632
rect 61838 -87646 61848 -87643
rect 61772 -87651 61848 -87646
rect 62134 -87650 62144 -87643
rect 62200 -87643 62500 -87612
rect 62200 -87650 62210 -87643
rect 62134 -87655 62210 -87650
rect 62490 -87646 62500 -87643
rect 62556 -87632 62840 -87606
rect 62934 -87622 63200 -86518
rect 63294 -87612 63560 -86508
rect 63654 -86500 63664 -86498
rect 63654 -86506 64364 -86500
rect 63654 -86508 63922 -86506
rect 63978 -86508 64276 -86506
rect 64332 -86508 64364 -86506
rect 63654 -87612 63910 -86508
rect 63294 -87622 63570 -87612
rect 62934 -87632 63210 -87622
rect 62556 -87643 62850 -87632
rect 62556 -87646 62566 -87643
rect 62490 -87651 62566 -87646
rect 62840 -87650 62850 -87643
rect 62906 -87643 63210 -87632
rect 62906 -87650 62916 -87643
rect 62840 -87655 62916 -87650
rect 63200 -87648 63210 -87643
rect 63266 -87643 63570 -87622
rect 63266 -87648 63276 -87643
rect 63200 -87653 63276 -87648
rect 63560 -87650 63570 -87643
rect 63626 -87622 63910 -87612
rect 64004 -87622 64270 -86508
rect 64364 -87622 64374 -86508
rect 68118 -87170 84140 -86520
rect 68118 -87172 68376 -87170
rect 77668 -87172 84140 -87170
rect 63626 -87643 63922 -87622
rect 63626 -87650 63636 -87643
rect 63912 -87644 63922 -87643
rect 63978 -87643 64276 -87622
rect 63978 -87644 63988 -87643
rect 63912 -87649 63988 -87644
rect 64266 -87644 64276 -87643
rect 64332 -87643 64364 -87622
rect 66300 -87632 67346 -87588
rect 66300 -87634 67028 -87632
rect 64332 -87644 64342 -87643
rect 64266 -87649 64342 -87644
rect 63560 -87655 63636 -87650
rect 66300 -87788 66316 -87634
rect 66372 -87788 66674 -87634
rect 66730 -87786 67028 -87634
rect 67084 -87786 67346 -87632
rect 66730 -87788 67346 -87786
rect 66300 -88060 67346 -87788
rect 68254 -87867 68314 -87858
rect 68610 -87863 68670 -87852
rect 66300 -88214 66324 -88060
rect 66380 -88062 67346 -88060
rect 66380 -88070 67038 -88062
rect 66380 -88214 66702 -88070
rect 66300 -88224 66702 -88214
rect 66758 -88216 67038 -88070
rect 67094 -88216 67346 -88062
rect 66758 -88224 67346 -88216
rect 66300 -88466 67346 -88224
rect 66300 -88620 66318 -88466
rect 66374 -88468 67346 -88466
rect 66374 -88472 67032 -88468
rect 66374 -88620 66674 -88472
rect 66300 -88626 66674 -88620
rect 66730 -88622 67032 -88472
rect 67088 -88622 67346 -88468
rect 66730 -88626 67346 -88622
rect 66300 -88880 67346 -88626
rect 66300 -89034 66318 -88880
rect 66374 -89034 66670 -88880
rect 66726 -89034 67032 -88880
rect 67088 -89034 67346 -88880
rect 68250 -87872 68328 -87867
rect 68250 -89024 68260 -87872
rect 68318 -89024 68328 -87872
rect 68430 -87868 68508 -87863
rect 68430 -87882 68440 -87868
rect 68498 -87882 68508 -87868
rect 68610 -87868 68696 -87863
rect 68426 -89014 68436 -87882
rect 68504 -89014 68514 -87882
rect 68250 -89029 68328 -89024
rect 68430 -89020 68440 -89014
rect 68498 -89020 68508 -89014
rect 68430 -89025 68508 -89020
rect 68610 -89020 68628 -87868
rect 68686 -89020 68696 -87868
rect 68968 -87867 69028 -87848
rect 68792 -87874 68870 -87869
rect 68792 -87890 68802 -87874
rect 68860 -87890 68870 -87874
rect 68968 -87872 69046 -87867
rect 69324 -87869 69384 -87852
rect 69682 -87867 69742 -87858
rect 68610 -89025 68696 -89020
rect 68788 -89022 68798 -87890
rect 68866 -89022 68876 -87890
rect 66300 -89068 67346 -89034
rect 54845 -90930 55821 -89292
rect 68254 -89295 68314 -89029
rect 68610 -89285 68670 -89025
rect 68792 -89026 68802 -89022
rect 68860 -89026 68870 -89022
rect 68792 -89031 68870 -89026
rect 68968 -89024 68978 -87872
rect 69036 -89024 69046 -87872
rect 69150 -87874 69228 -87869
rect 69150 -87890 69160 -87874
rect 69138 -89022 69148 -87890
rect 68968 -89029 69046 -89024
rect 69150 -89026 69160 -89022
rect 69218 -89026 69228 -87874
rect 68434 -89294 68512 -89289
rect 68254 -89300 68336 -89295
rect 56532 -89338 56612 -89333
rect 56532 -89346 56542 -89338
rect 56602 -89346 56612 -89338
rect 56890 -89336 56970 -89331
rect 58672 -89334 58752 -89329
rect 59736 -89330 59816 -89325
rect 56890 -89342 56900 -89336
rect 56960 -89342 56970 -89336
rect 57244 -89342 57324 -89337
rect 56524 -90468 56534 -89346
rect 56610 -90468 56620 -89346
rect 56884 -90464 56894 -89342
rect 56970 -90464 56980 -89342
rect 57244 -89352 57254 -89342
rect 57314 -89352 57324 -89342
rect 57598 -89348 57678 -89343
rect 57598 -89352 57608 -89348
rect 57668 -89352 57678 -89348
rect 57954 -89344 58034 -89339
rect 57954 -89350 57964 -89344
rect 58024 -89350 58034 -89344
rect 58312 -89340 58392 -89335
rect 58672 -89338 58682 -89334
rect 58742 -89338 58752 -89334
rect 59378 -89338 59458 -89333
rect 59736 -89334 59746 -89330
rect 59806 -89334 59816 -89330
rect 61670 -89334 61750 -89329
rect 58312 -89348 58322 -89340
rect 58382 -89348 58392 -89340
rect 56532 -90472 56542 -90468
rect 56602 -90472 56612 -90468
rect 56532 -90477 56612 -90472
rect 56890 -90470 56900 -90464
rect 56960 -90470 56970 -90464
rect 56890 -90475 56970 -90470
rect 57240 -90474 57250 -89352
rect 57326 -90474 57336 -89352
rect 57590 -90474 57600 -89352
rect 57676 -90474 57686 -89352
rect 57946 -90472 57956 -89350
rect 58032 -90472 58042 -89350
rect 58302 -90470 58312 -89348
rect 58388 -90470 58398 -89348
rect 58664 -90460 58674 -89338
rect 58750 -90460 58760 -89338
rect 59378 -89340 59388 -89338
rect 59448 -89340 59458 -89338
rect 59018 -89346 59098 -89341
rect 59018 -89350 59028 -89346
rect 59088 -89350 59098 -89346
rect 58672 -90468 58682 -90460
rect 58742 -90468 58752 -90460
rect 57244 -90476 57254 -90474
rect 57314 -90476 57324 -90474
rect 57244 -90481 57324 -90476
rect 57598 -90482 57608 -90474
rect 57668 -90482 57678 -90474
rect 57598 -90487 57678 -90482
rect 57954 -90478 57964 -90472
rect 58024 -90478 58034 -90472
rect 57954 -90483 58034 -90478
rect 58312 -90474 58322 -90470
rect 58382 -90474 58392 -90470
rect 58672 -90473 58752 -90468
rect 59014 -90472 59024 -89350
rect 59100 -90472 59110 -89350
rect 59376 -90462 59386 -89340
rect 59462 -90462 59472 -89340
rect 59726 -90456 59736 -89334
rect 59812 -90456 59822 -89334
rect 60964 -89340 61044 -89335
rect 60964 -89342 60974 -89340
rect 61034 -89342 61044 -89340
rect 61312 -89342 61392 -89337
rect 61670 -89338 61680 -89334
rect 61740 -89338 61750 -89334
rect 60954 -89770 60964 -89342
rect 59378 -90472 59388 -90462
rect 59448 -90472 59458 -90462
rect 59736 -90464 59746 -90456
rect 59806 -90464 59816 -90456
rect 59736 -90469 59816 -90464
rect 60756 -90464 60964 -89770
rect 61040 -89770 61050 -89342
rect 61312 -89352 61322 -89342
rect 61382 -89352 61392 -89342
rect 61308 -89770 61318 -89352
rect 61040 -90464 61318 -89770
rect 58312 -90479 58392 -90474
rect 59018 -90480 59028 -90472
rect 59088 -90480 59098 -90472
rect 59378 -90477 59458 -90472
rect 60756 -90474 60974 -90464
rect 61034 -90474 61318 -90464
rect 61394 -89770 61404 -89352
rect 61666 -89770 61676 -89338
rect 61394 -90460 61676 -89770
rect 61752 -89770 61762 -89338
rect 62032 -89344 62112 -89339
rect 63096 -89340 63176 -89335
rect 62032 -89348 62042 -89344
rect 62102 -89348 62112 -89344
rect 62386 -89348 62466 -89343
rect 62026 -89770 62036 -89348
rect 61752 -90460 62036 -89770
rect 61394 -90468 61680 -90460
rect 61740 -90468 62036 -90460
rect 61394 -90470 62036 -90468
rect 62112 -89770 62122 -89348
rect 62386 -89354 62396 -89348
rect 62456 -89354 62466 -89348
rect 62742 -89348 62822 -89343
rect 63096 -89346 63106 -89340
rect 63166 -89346 63176 -89340
rect 63816 -89344 63896 -89339
rect 63816 -89346 63826 -89344
rect 63886 -89346 63896 -89344
rect 62742 -89352 62752 -89348
rect 62812 -89352 62822 -89348
rect 62382 -89770 62392 -89354
rect 62112 -90470 62392 -89770
rect 61394 -90474 62042 -90470
rect 60756 -90476 61322 -90474
rect 61382 -90476 62042 -90474
rect 59018 -90485 59098 -90480
rect 60756 -90478 62042 -90476
rect 62102 -90476 62392 -90470
rect 62468 -89770 62478 -89354
rect 62732 -89770 62742 -89352
rect 62468 -90474 62742 -89770
rect 62818 -89770 62828 -89352
rect 63094 -89770 63104 -89346
rect 62818 -90468 63104 -89770
rect 63180 -89770 63190 -89346
rect 63456 -89352 63536 -89347
rect 63456 -89360 63466 -89352
rect 63526 -89360 63536 -89352
rect 63448 -89770 63458 -89360
rect 63180 -90468 63458 -89770
rect 62818 -90474 63106 -90468
rect 63166 -90474 63458 -90468
rect 62468 -90476 62752 -90474
rect 62102 -90478 62396 -90476
rect 60756 -90482 62396 -90478
rect 62456 -90482 62752 -90476
rect 62812 -90482 63458 -90474
rect 63534 -89770 63544 -89360
rect 63806 -89770 63816 -89346
rect 63534 -90468 63816 -89770
rect 63892 -89770 63902 -89346
rect 64172 -89348 64252 -89343
rect 64172 -89352 64182 -89348
rect 64242 -89352 64252 -89348
rect 64166 -89770 64176 -89352
rect 63892 -90468 64176 -89770
rect 63534 -90478 63826 -90468
rect 63886 -90474 64176 -90468
rect 64252 -89770 64262 -89352
rect 64252 -90474 66766 -89770
rect 63886 -90478 64182 -90474
rect 63534 -90482 64182 -90478
rect 64242 -90482 66766 -90474
rect 60756 -90486 63466 -90482
rect 63526 -90486 66766 -90482
rect 60756 -90530 66766 -90486
rect 68254 -90452 68268 -89300
rect 68326 -90452 68336 -89300
rect 68434 -89308 68444 -89294
rect 68502 -89308 68512 -89294
rect 68610 -89290 68690 -89285
rect 68430 -90440 68440 -89308
rect 68508 -90440 68518 -89308
rect 68434 -90446 68444 -90440
rect 68502 -90446 68512 -90440
rect 68434 -90451 68512 -90446
rect 68610 -90442 68622 -89290
rect 68680 -90442 68690 -89290
rect 68790 -89296 68868 -89291
rect 68790 -89308 68800 -89296
rect 68858 -89308 68868 -89296
rect 68968 -89293 69028 -89029
rect 69150 -89031 69228 -89026
rect 69324 -87874 69406 -87869
rect 69324 -89026 69338 -87874
rect 69396 -89026 69406 -87874
rect 69502 -87872 69580 -87867
rect 69502 -87892 69512 -87872
rect 69570 -87892 69580 -87872
rect 69682 -87872 69760 -87867
rect 69496 -89024 69506 -87892
rect 69574 -89024 69584 -87892
rect 69682 -89024 69692 -87872
rect 69750 -89024 69760 -87872
rect 69856 -87874 69934 -87869
rect 69856 -87888 69866 -87874
rect 69924 -87888 69934 -87874
rect 70036 -87873 70096 -87852
rect 70394 -87867 70454 -87858
rect 70390 -87872 70468 -87867
rect 70036 -87878 70116 -87873
rect 69850 -89020 69860 -87888
rect 69928 -89020 69938 -87888
rect 69324 -89031 69406 -89026
rect 69502 -89029 69580 -89024
rect 69682 -89029 69760 -89024
rect 69856 -89026 69866 -89020
rect 69924 -89026 69934 -89020
rect 68968 -89298 69048 -89293
rect 68786 -90440 68796 -89308
rect 68864 -90440 68874 -89308
rect 68610 -90447 68690 -90442
rect 68254 -90457 68336 -90452
rect 68254 -90930 68314 -90457
rect 68610 -90930 68670 -90447
rect 68790 -90448 68800 -90440
rect 68858 -90448 68868 -90440
rect 68790 -90453 68868 -90448
rect 68968 -90450 68980 -89298
rect 69038 -90450 69048 -89298
rect 69146 -89294 69224 -89289
rect 69324 -89293 69384 -89031
rect 69498 -89292 69576 -89287
rect 69682 -89289 69742 -89029
rect 69856 -89031 69934 -89026
rect 70036 -89030 70048 -87878
rect 70106 -89030 70116 -87878
rect 70212 -87880 70290 -87875
rect 70212 -87894 70222 -87880
rect 70202 -89026 70212 -87894
rect 70036 -89035 70116 -89030
rect 70212 -89032 70222 -89026
rect 70280 -89032 70290 -87880
rect 70390 -89024 70400 -87872
rect 70458 -89024 70468 -87872
rect 70750 -87873 70810 -87868
rect 71100 -87871 71160 -87858
rect 70572 -87878 70650 -87873
rect 70572 -87890 70582 -87878
rect 70640 -87890 70650 -87878
rect 70746 -87878 70824 -87873
rect 70564 -89022 70574 -87890
rect 70642 -89022 70652 -87890
rect 70390 -89029 70468 -89024
rect 70036 -89289 70096 -89035
rect 70212 -89037 70290 -89032
rect 69146 -89308 69156 -89294
rect 69214 -89308 69224 -89294
rect 69322 -89298 69400 -89293
rect 69140 -90440 69150 -89308
rect 69218 -90440 69228 -89308
rect 68968 -90455 69048 -90450
rect 69146 -90446 69156 -90440
rect 69214 -90446 69224 -90440
rect 69146 -90451 69224 -90446
rect 69322 -90450 69332 -89298
rect 69390 -90450 69400 -89298
rect 69498 -89310 69508 -89292
rect 69566 -89310 69576 -89292
rect 69678 -89294 69756 -89289
rect 69490 -90442 69500 -89310
rect 69568 -90442 69578 -89310
rect 69498 -90444 69508 -90442
rect 69566 -90444 69576 -90442
rect 69498 -90449 69576 -90444
rect 69678 -90446 69688 -89294
rect 69746 -90446 69756 -89294
rect 69854 -89298 69932 -89293
rect 69854 -89316 69864 -89298
rect 69922 -89316 69932 -89298
rect 70034 -89294 70112 -89289
rect 69322 -90455 69400 -90450
rect 69678 -90451 69756 -90446
rect 69846 -90448 69856 -89316
rect 69924 -90448 69934 -89316
rect 70034 -90446 70044 -89294
rect 70102 -90446 70112 -89294
rect 70216 -89292 70294 -89287
rect 70216 -89316 70226 -89292
rect 70284 -89316 70294 -89292
rect 70394 -89289 70454 -89029
rect 70572 -89030 70582 -89022
rect 70640 -89030 70650 -89022
rect 70572 -89035 70650 -89030
rect 70746 -89030 70756 -87878
rect 70814 -89030 70824 -87878
rect 70926 -87876 71004 -87871
rect 70926 -87894 70936 -87876
rect 70994 -87894 71004 -87876
rect 71100 -87876 71186 -87871
rect 70918 -89026 70928 -87894
rect 70996 -89026 71006 -87894
rect 70746 -89035 70824 -89030
rect 70926 -89028 70936 -89026
rect 70994 -89028 71004 -89026
rect 70926 -89033 71004 -89028
rect 71100 -89028 71118 -87876
rect 71176 -89028 71186 -87876
rect 71458 -87875 71518 -87852
rect 71814 -87871 71874 -87852
rect 74144 -87865 74204 -87846
rect 74500 -87861 74560 -87852
rect 74144 -87870 74224 -87865
rect 71282 -87882 71360 -87877
rect 71282 -87898 71292 -87882
rect 71350 -87898 71360 -87882
rect 71458 -87880 71540 -87875
rect 71100 -89033 71186 -89028
rect 71276 -89030 71286 -87898
rect 71354 -89030 71364 -87898
rect 70750 -89289 70810 -89035
rect 71100 -89283 71160 -89033
rect 71282 -89034 71292 -89030
rect 71350 -89034 71360 -89030
rect 71282 -89039 71360 -89034
rect 71458 -89032 71472 -87880
rect 71530 -89032 71540 -87880
rect 71636 -87880 71714 -87875
rect 71636 -87894 71646 -87880
rect 71704 -87894 71714 -87880
rect 71814 -87876 71892 -87871
rect 71634 -89026 71644 -87894
rect 71712 -89026 71722 -87894
rect 71458 -89037 71540 -89032
rect 71636 -89032 71646 -89026
rect 71704 -89032 71714 -89026
rect 71636 -89037 71714 -89032
rect 71814 -89028 71824 -87876
rect 71882 -89028 71892 -87876
rect 71814 -89033 71892 -89028
rect 74144 -89022 74156 -87870
rect 74214 -89022 74224 -87870
rect 74326 -87866 74404 -87861
rect 74326 -87880 74336 -87866
rect 74394 -87880 74404 -87866
rect 74500 -87866 74592 -87861
rect 74322 -89012 74332 -87880
rect 74400 -89012 74410 -87880
rect 74144 -89027 74224 -89022
rect 74326 -89018 74336 -89012
rect 74394 -89018 74404 -89012
rect 74326 -89023 74404 -89018
rect 74500 -89018 74524 -87866
rect 74582 -89018 74592 -87866
rect 74858 -87865 74918 -87852
rect 74688 -87872 74766 -87867
rect 74688 -87888 74698 -87872
rect 74756 -87888 74766 -87872
rect 74858 -87870 74942 -87865
rect 75214 -87867 75274 -87854
rect 75572 -87865 75632 -87854
rect 74500 -89023 74592 -89018
rect 74684 -89020 74694 -87888
rect 74762 -89020 74772 -87888
rect 71100 -89288 71180 -89283
rect 70394 -89294 70474 -89289
rect 69854 -90450 69864 -90448
rect 69922 -90450 69932 -90448
rect 68968 -90930 69028 -90455
rect 69324 -90930 69384 -90455
rect 69682 -90930 69742 -90451
rect 69854 -90455 69932 -90450
rect 70034 -90451 70112 -90446
rect 70210 -90448 70220 -89316
rect 70288 -90448 70298 -89316
rect 70394 -90446 70406 -89294
rect 70464 -90446 70474 -89294
rect 70568 -89294 70646 -89289
rect 70568 -89314 70578 -89294
rect 70636 -89314 70646 -89294
rect 70746 -89294 70824 -89289
rect 70560 -90446 70570 -89314
rect 70638 -90446 70648 -89314
rect 70746 -90446 70756 -89294
rect 70814 -90446 70824 -89294
rect 70924 -89294 71002 -89289
rect 70924 -89312 70934 -89294
rect 70992 -89312 71002 -89294
rect 70916 -90444 70926 -89312
rect 70994 -90444 71004 -89312
rect 71100 -90440 71112 -89288
rect 71170 -90440 71180 -89288
rect 71284 -89298 71362 -89293
rect 71284 -89316 71294 -89298
rect 71352 -89316 71362 -89298
rect 71458 -89295 71518 -89037
rect 71636 -89294 71714 -89289
rect 71458 -89300 71540 -89295
rect 70216 -90449 70294 -90448
rect 70394 -90451 70474 -90446
rect 70568 -90451 70646 -90446
rect 70746 -90451 70824 -90446
rect 70924 -90446 70934 -90444
rect 70992 -90446 71002 -90444
rect 70924 -90451 71002 -90446
rect 71100 -90445 71180 -90440
rect 70036 -90930 70096 -90451
rect 70394 -90930 70454 -90451
rect 70750 -90930 70810 -90451
rect 71100 -90930 71160 -90445
rect 71276 -90448 71286 -89316
rect 71354 -90448 71364 -89316
rect 71284 -90450 71294 -90448
rect 71352 -90450 71362 -90448
rect 71284 -90455 71362 -90450
rect 71458 -90452 71472 -89300
rect 71530 -90452 71540 -89300
rect 71636 -89316 71646 -89294
rect 71624 -90448 71634 -89316
rect 71704 -90446 71714 -89294
rect 71702 -90448 71714 -90446
rect 71636 -90451 71714 -90448
rect 71814 -89293 71874 -89033
rect 74144 -89293 74204 -89027
rect 74500 -89283 74560 -89023
rect 74688 -89024 74698 -89020
rect 74756 -89024 74766 -89020
rect 74688 -89029 74766 -89024
rect 74858 -89022 74874 -87870
rect 74932 -89022 74942 -87870
rect 75046 -87872 75124 -87867
rect 75046 -87888 75056 -87872
rect 75034 -89020 75044 -87888
rect 74858 -89027 74942 -89022
rect 75046 -89024 75056 -89020
rect 75114 -89024 75124 -87872
rect 74330 -89292 74408 -89287
rect 71814 -89298 71894 -89293
rect 71814 -90450 71826 -89298
rect 71884 -90450 71894 -89298
rect 71458 -90457 71540 -90452
rect 71814 -90455 71894 -90450
rect 74144 -89298 74232 -89293
rect 74144 -90450 74164 -89298
rect 74222 -90450 74232 -89298
rect 74330 -89306 74340 -89292
rect 74398 -89306 74408 -89292
rect 74500 -89288 74586 -89283
rect 74326 -90438 74336 -89306
rect 74404 -90438 74414 -89306
rect 74330 -90444 74340 -90438
rect 74398 -90444 74408 -90438
rect 74330 -90449 74408 -90444
rect 74500 -90440 74518 -89288
rect 74576 -90440 74586 -89288
rect 74686 -89294 74764 -89289
rect 74686 -89306 74696 -89294
rect 74754 -89306 74764 -89294
rect 74858 -89291 74918 -89027
rect 75046 -89029 75124 -89024
rect 75214 -87872 75302 -87867
rect 75214 -89024 75234 -87872
rect 75292 -89024 75302 -87872
rect 75398 -87870 75476 -87865
rect 75398 -87890 75408 -87870
rect 75466 -87890 75476 -87870
rect 75572 -87870 75656 -87865
rect 75392 -89022 75402 -87890
rect 75470 -89022 75480 -87890
rect 75572 -89022 75588 -87870
rect 75646 -89022 75656 -87870
rect 75752 -87872 75830 -87867
rect 75752 -87886 75762 -87872
rect 75820 -87886 75830 -87872
rect 75926 -87871 75986 -87854
rect 76284 -87865 76344 -87840
rect 76284 -87870 76364 -87865
rect 75926 -87876 76012 -87871
rect 75746 -89018 75756 -87886
rect 75824 -89018 75834 -87886
rect 75214 -89029 75302 -89024
rect 75398 -89027 75476 -89022
rect 75572 -89027 75656 -89022
rect 75752 -89024 75762 -89018
rect 75820 -89024 75830 -89018
rect 74858 -89296 74944 -89291
rect 74682 -90438 74692 -89306
rect 74760 -90438 74770 -89306
rect 74500 -90445 74586 -90440
rect 74144 -90455 74232 -90450
rect 71458 -90930 71518 -90457
rect 71814 -90930 71874 -90455
rect 74144 -90930 74204 -90455
rect 74500 -90930 74560 -90445
rect 74686 -90446 74696 -90438
rect 74754 -90446 74764 -90438
rect 74686 -90451 74764 -90446
rect 74858 -90448 74876 -89296
rect 74934 -90448 74944 -89296
rect 75042 -89292 75120 -89287
rect 75042 -89306 75052 -89292
rect 75110 -89306 75120 -89292
rect 75214 -89291 75274 -89029
rect 75394 -89290 75472 -89285
rect 75214 -89296 75296 -89291
rect 75036 -90438 75046 -89306
rect 75114 -90438 75124 -89306
rect 74858 -90453 74944 -90448
rect 75042 -90444 75052 -90438
rect 75110 -90444 75120 -90438
rect 75042 -90449 75120 -90444
rect 75214 -90448 75228 -89296
rect 75286 -90448 75296 -89296
rect 75394 -89308 75404 -89290
rect 75462 -89308 75472 -89290
rect 75572 -89287 75632 -89027
rect 75752 -89029 75830 -89024
rect 75926 -89028 75944 -87876
rect 76002 -89028 76012 -87876
rect 76108 -87878 76186 -87873
rect 76108 -87892 76118 -87878
rect 76098 -89024 76108 -87892
rect 75926 -89033 76012 -89028
rect 76108 -89030 76118 -89024
rect 76176 -89030 76186 -87878
rect 75926 -89287 75986 -89033
rect 76108 -89035 76186 -89030
rect 76284 -89022 76296 -87870
rect 76354 -89022 76364 -87870
rect 76640 -87871 76700 -87854
rect 76990 -87869 77050 -87854
rect 76468 -87876 76546 -87871
rect 76468 -87888 76478 -87876
rect 76536 -87888 76546 -87876
rect 76640 -87876 76720 -87871
rect 76460 -89020 76470 -87888
rect 76538 -89020 76548 -87888
rect 76284 -89027 76364 -89022
rect 75572 -89292 75652 -89287
rect 75386 -90440 75396 -89308
rect 75464 -90440 75474 -89308
rect 75394 -90442 75404 -90440
rect 75462 -90442 75472 -90440
rect 75394 -90447 75472 -90442
rect 75572 -90444 75584 -89292
rect 75642 -90444 75652 -89292
rect 75750 -89296 75828 -89291
rect 75750 -89314 75760 -89296
rect 75818 -89314 75828 -89296
rect 75926 -89292 76008 -89287
rect 75214 -90453 75296 -90448
rect 75572 -90449 75652 -90444
rect 75742 -90446 75752 -89314
rect 75820 -90446 75830 -89314
rect 75926 -90444 75940 -89292
rect 75998 -90444 76008 -89292
rect 76112 -89290 76190 -89285
rect 76112 -89314 76122 -89290
rect 76180 -89314 76190 -89290
rect 76284 -89287 76344 -89027
rect 76468 -89028 76478 -89020
rect 76536 -89028 76546 -89020
rect 76468 -89033 76546 -89028
rect 76640 -89028 76652 -87876
rect 76710 -89028 76720 -87876
rect 76822 -87874 76900 -87869
rect 76822 -87892 76832 -87874
rect 76890 -87892 76900 -87874
rect 76990 -87874 77082 -87869
rect 76814 -89024 76824 -87892
rect 76892 -89024 76902 -87892
rect 76640 -89033 76720 -89028
rect 76822 -89026 76832 -89024
rect 76890 -89026 76900 -89024
rect 76822 -89031 76900 -89026
rect 76990 -89026 77014 -87874
rect 77072 -89026 77082 -87874
rect 77348 -87873 77408 -87854
rect 77704 -87869 77764 -87848
rect 80274 -87859 80334 -87848
rect 80630 -87855 80690 -87854
rect 80260 -87864 80338 -87859
rect 77178 -87880 77256 -87875
rect 77178 -87896 77188 -87880
rect 77246 -87896 77256 -87880
rect 77348 -87878 77436 -87873
rect 76990 -89031 77082 -89026
rect 77172 -89028 77182 -87896
rect 77250 -89028 77260 -87896
rect 76640 -89287 76700 -89033
rect 76990 -89281 77050 -89031
rect 77178 -89032 77188 -89028
rect 77246 -89032 77256 -89028
rect 77178 -89037 77256 -89032
rect 77348 -89030 77368 -87878
rect 77426 -89030 77436 -87878
rect 77532 -87878 77610 -87873
rect 77532 -87892 77542 -87878
rect 77600 -87892 77610 -87878
rect 77704 -87874 77788 -87869
rect 77530 -89024 77540 -87892
rect 77608 -89024 77618 -87892
rect 77348 -89035 77436 -89030
rect 77532 -89030 77542 -89024
rect 77600 -89030 77610 -89024
rect 77532 -89035 77610 -89030
rect 77704 -89026 77720 -87874
rect 77778 -89026 77788 -87874
rect 80260 -89016 80270 -87864
rect 80328 -89016 80338 -87864
rect 80440 -87860 80518 -87855
rect 80440 -87874 80450 -87860
rect 80508 -87874 80518 -87860
rect 80628 -87860 80706 -87855
rect 80988 -87859 81048 -87848
rect 80436 -89006 80446 -87874
rect 80514 -89006 80524 -87874
rect 80260 -89021 80338 -89016
rect 80440 -89012 80450 -89006
rect 80508 -89012 80518 -89006
rect 80440 -89017 80518 -89012
rect 80628 -89012 80638 -87860
rect 80696 -89012 80706 -87860
rect 80802 -87866 80880 -87861
rect 80802 -87882 80812 -87866
rect 80870 -87882 80880 -87866
rect 80978 -87864 81056 -87859
rect 81344 -87861 81404 -87848
rect 81702 -87859 81762 -87848
rect 80628 -89017 80706 -89012
rect 80798 -89014 80808 -87882
rect 80876 -89014 80886 -87882
rect 77704 -89031 77788 -89026
rect 76990 -89286 77076 -89281
rect 76284 -89292 76370 -89287
rect 75750 -90448 75760 -90446
rect 75818 -90448 75828 -90446
rect 74858 -90930 74918 -90453
rect 75214 -90930 75274 -90453
rect 75572 -90930 75632 -90449
rect 75750 -90453 75828 -90448
rect 75926 -90449 76008 -90444
rect 76106 -90446 76116 -89314
rect 76184 -90446 76194 -89314
rect 76284 -90444 76302 -89292
rect 76360 -90444 76370 -89292
rect 76464 -89292 76542 -89287
rect 76464 -89312 76474 -89292
rect 76532 -89312 76542 -89292
rect 76640 -89292 76720 -89287
rect 76456 -90444 76466 -89312
rect 76534 -90444 76544 -89312
rect 76640 -90444 76652 -89292
rect 76710 -90444 76720 -89292
rect 76820 -89292 76898 -89287
rect 76820 -89310 76830 -89292
rect 76888 -89310 76898 -89292
rect 76812 -90442 76822 -89310
rect 76890 -90442 76900 -89310
rect 76990 -90438 77008 -89286
rect 77066 -90438 77076 -89286
rect 77180 -89296 77258 -89291
rect 77180 -89314 77190 -89296
rect 77248 -89314 77258 -89296
rect 77348 -89293 77408 -89035
rect 77532 -89292 77610 -89287
rect 77348 -89298 77436 -89293
rect 76112 -90447 76190 -90446
rect 76284 -90449 76370 -90444
rect 76464 -90449 76542 -90444
rect 76640 -90449 76720 -90444
rect 76820 -90444 76830 -90442
rect 76888 -90444 76898 -90442
rect 76820 -90449 76898 -90444
rect 76990 -90443 77076 -90438
rect 75926 -90930 75986 -90449
rect 76284 -90930 76344 -90449
rect 76640 -90930 76700 -90449
rect 76990 -90930 77050 -90443
rect 77172 -90446 77182 -89314
rect 77250 -90446 77260 -89314
rect 77180 -90448 77190 -90446
rect 77248 -90448 77258 -90446
rect 77180 -90453 77258 -90448
rect 77348 -90450 77368 -89298
rect 77426 -90450 77436 -89298
rect 77532 -89314 77542 -89292
rect 77520 -90446 77530 -89314
rect 77600 -90444 77610 -89292
rect 77598 -90446 77610 -90444
rect 77532 -90449 77610 -90446
rect 77704 -89291 77764 -89031
rect 80274 -89287 80334 -89021
rect 80630 -89277 80690 -89017
rect 80802 -89018 80812 -89014
rect 80870 -89018 80880 -89014
rect 80802 -89023 80880 -89018
rect 80978 -89016 80988 -87864
rect 81046 -89016 81056 -87864
rect 81160 -87866 81238 -87861
rect 81160 -87882 81170 -87866
rect 81148 -89014 81158 -87882
rect 80978 -89021 81056 -89016
rect 81160 -89018 81170 -89014
rect 81228 -89018 81238 -87866
rect 80444 -89286 80522 -89281
rect 77704 -89296 77790 -89291
rect 77704 -90448 77722 -89296
rect 77780 -90448 77790 -89296
rect 77348 -90455 77436 -90450
rect 77704 -90453 77790 -90448
rect 80268 -89292 80346 -89287
rect 80268 -90444 80278 -89292
rect 80336 -90444 80346 -89292
rect 80444 -89300 80454 -89286
rect 80512 -89300 80522 -89286
rect 80622 -89282 80700 -89277
rect 80440 -90432 80450 -89300
rect 80518 -90432 80528 -89300
rect 80444 -90438 80454 -90432
rect 80512 -90438 80522 -90432
rect 80444 -90443 80522 -90438
rect 80622 -90434 80632 -89282
rect 80690 -90434 80700 -89282
rect 80800 -89288 80878 -89283
rect 80988 -89285 81048 -89021
rect 81160 -89023 81238 -89018
rect 81338 -87866 81416 -87861
rect 81338 -89018 81348 -87866
rect 81406 -89018 81416 -87866
rect 81512 -87864 81590 -87859
rect 81512 -87884 81522 -87864
rect 81580 -87884 81590 -87864
rect 81692 -87864 81770 -87859
rect 81506 -89016 81516 -87884
rect 81584 -89016 81594 -87884
rect 81692 -89016 81702 -87864
rect 81760 -89016 81770 -87864
rect 81866 -87866 81944 -87861
rect 82056 -87865 82116 -87848
rect 82414 -87859 82474 -87854
rect 82400 -87864 82478 -87859
rect 81866 -87880 81876 -87866
rect 81934 -87880 81944 -87866
rect 82048 -87870 82126 -87865
rect 81860 -89012 81870 -87880
rect 81938 -89012 81948 -87880
rect 81338 -89023 81416 -89018
rect 81512 -89021 81590 -89016
rect 81692 -89021 81770 -89016
rect 81866 -89018 81876 -89012
rect 81934 -89018 81944 -89012
rect 80800 -89300 80810 -89288
rect 80868 -89300 80878 -89288
rect 80980 -89290 81058 -89285
rect 80796 -90432 80806 -89300
rect 80874 -90432 80884 -89300
rect 80622 -90439 80700 -90434
rect 80268 -90449 80346 -90444
rect 77348 -90930 77408 -90455
rect 77704 -90930 77764 -90453
rect 80274 -90930 80334 -90449
rect 80630 -90930 80690 -90439
rect 80800 -90440 80810 -90432
rect 80868 -90440 80878 -90432
rect 80800 -90445 80878 -90440
rect 80980 -90442 80990 -89290
rect 81048 -90442 81058 -89290
rect 81156 -89286 81234 -89281
rect 81344 -89285 81404 -89023
rect 81508 -89284 81586 -89279
rect 81702 -89281 81762 -89021
rect 81866 -89023 81944 -89018
rect 82048 -89022 82058 -87870
rect 82116 -89022 82126 -87870
rect 82222 -87872 82300 -87867
rect 82222 -87886 82232 -87872
rect 82212 -89018 82222 -87886
rect 82048 -89027 82126 -89022
rect 82222 -89024 82232 -89018
rect 82290 -89024 82300 -87872
rect 82400 -89016 82410 -87864
rect 82468 -89016 82478 -87864
rect 82770 -87865 82830 -87840
rect 83120 -87863 83180 -87848
rect 82582 -87870 82660 -87865
rect 82582 -87882 82592 -87870
rect 82650 -87882 82660 -87870
rect 82756 -87870 82834 -87865
rect 82574 -89014 82584 -87882
rect 82652 -89014 82662 -87882
rect 82400 -89021 82478 -89016
rect 82056 -89281 82116 -89027
rect 82222 -89029 82300 -89024
rect 81156 -89300 81166 -89286
rect 81224 -89300 81234 -89286
rect 81332 -89290 81410 -89285
rect 81150 -90432 81160 -89300
rect 81228 -90432 81238 -89300
rect 80980 -90447 81058 -90442
rect 81156 -90438 81166 -90432
rect 81224 -90438 81234 -90432
rect 81156 -90443 81234 -90438
rect 81332 -90442 81342 -89290
rect 81400 -90442 81410 -89290
rect 81508 -89302 81518 -89284
rect 81576 -89302 81586 -89284
rect 81688 -89286 81766 -89281
rect 81500 -90434 81510 -89302
rect 81578 -90434 81588 -89302
rect 81508 -90436 81518 -90434
rect 81576 -90436 81586 -90434
rect 81508 -90441 81586 -90436
rect 81688 -90438 81698 -89286
rect 81756 -90438 81766 -89286
rect 81864 -89290 81942 -89285
rect 81864 -89308 81874 -89290
rect 81932 -89308 81942 -89290
rect 82044 -89286 82122 -89281
rect 81332 -90447 81410 -90442
rect 81688 -90443 81766 -90438
rect 81856 -90440 81866 -89308
rect 81934 -90440 81944 -89308
rect 82044 -90438 82054 -89286
rect 82112 -90438 82122 -89286
rect 82226 -89284 82304 -89279
rect 82414 -89281 82474 -89021
rect 82582 -89022 82592 -89014
rect 82650 -89022 82660 -89014
rect 82582 -89027 82660 -89022
rect 82756 -89022 82766 -87870
rect 82824 -89022 82834 -87870
rect 82936 -87868 83014 -87863
rect 82936 -87886 82946 -87868
rect 83004 -87886 83014 -87868
rect 83118 -87868 83196 -87863
rect 83478 -87867 83538 -87840
rect 83834 -87863 83894 -87848
rect 82928 -89018 82938 -87886
rect 83006 -89018 83016 -87886
rect 82756 -89027 82834 -89022
rect 82936 -89020 82946 -89018
rect 83004 -89020 83014 -89018
rect 82936 -89025 83014 -89020
rect 83118 -89020 83128 -87868
rect 83186 -89020 83196 -87868
rect 83292 -87874 83370 -87869
rect 83292 -87890 83302 -87874
rect 83360 -87890 83370 -87874
rect 83472 -87872 83550 -87867
rect 83118 -89025 83196 -89020
rect 83286 -89022 83296 -87890
rect 83364 -89022 83374 -87890
rect 82770 -89281 82830 -89027
rect 83120 -89275 83180 -89025
rect 83292 -89026 83302 -89022
rect 83360 -89026 83370 -89022
rect 83292 -89031 83370 -89026
rect 83472 -89024 83482 -87872
rect 83540 -89024 83550 -87872
rect 83646 -87872 83724 -87867
rect 83646 -87886 83656 -87872
rect 83714 -87886 83724 -87872
rect 83824 -87868 83902 -87863
rect 83644 -89018 83654 -87886
rect 83722 -89018 83732 -87886
rect 83472 -89029 83550 -89024
rect 83646 -89024 83656 -89018
rect 83714 -89024 83724 -89018
rect 83646 -89029 83724 -89024
rect 83824 -89020 83834 -87868
rect 83892 -89020 83902 -87868
rect 83824 -89025 83902 -89020
rect 83112 -89280 83190 -89275
rect 82226 -89308 82236 -89284
rect 82294 -89308 82304 -89284
rect 82406 -89286 82484 -89281
rect 81864 -90442 81874 -90440
rect 81932 -90442 81942 -90440
rect 80988 -90930 81048 -90447
rect 81344 -90930 81404 -90447
rect 81702 -90930 81762 -90443
rect 81864 -90447 81942 -90442
rect 82044 -90443 82122 -90438
rect 82220 -90440 82230 -89308
rect 82298 -90440 82308 -89308
rect 82406 -90438 82416 -89286
rect 82474 -90438 82484 -89286
rect 82578 -89286 82656 -89281
rect 82578 -89306 82588 -89286
rect 82646 -89306 82656 -89286
rect 82756 -89286 82834 -89281
rect 82570 -90438 82580 -89306
rect 82648 -90438 82658 -89306
rect 82756 -90438 82766 -89286
rect 82824 -90438 82834 -89286
rect 82934 -89286 83012 -89281
rect 82934 -89304 82944 -89286
rect 83002 -89304 83012 -89286
rect 82926 -90436 82936 -89304
rect 83004 -90436 83014 -89304
rect 83112 -90432 83122 -89280
rect 83180 -90432 83190 -89280
rect 83294 -89290 83372 -89285
rect 83478 -89287 83538 -89029
rect 83646 -89286 83724 -89281
rect 83834 -89285 83894 -89025
rect 83294 -89308 83304 -89290
rect 83362 -89308 83372 -89290
rect 83472 -89292 83550 -89287
rect 82226 -90441 82304 -90440
rect 82406 -90443 82484 -90438
rect 82578 -90443 82656 -90438
rect 82756 -90443 82834 -90438
rect 82934 -90438 82944 -90436
rect 83002 -90438 83012 -90436
rect 83112 -90437 83190 -90432
rect 82934 -90443 83012 -90438
rect 82056 -90930 82116 -90443
rect 82414 -90930 82474 -90443
rect 82770 -90930 82830 -90443
rect 83120 -90930 83180 -90437
rect 83286 -90440 83296 -89308
rect 83364 -90440 83374 -89308
rect 83294 -90442 83304 -90440
rect 83362 -90442 83372 -90440
rect 83294 -90447 83372 -90442
rect 83472 -90444 83482 -89292
rect 83540 -90444 83550 -89292
rect 83646 -89308 83656 -89286
rect 83634 -90440 83644 -89308
rect 83714 -90438 83724 -89286
rect 83712 -90440 83724 -90438
rect 83646 -90443 83724 -90440
rect 83826 -89290 83904 -89285
rect 83826 -90442 83836 -89290
rect 83894 -90442 83904 -89290
rect 83472 -90449 83550 -90444
rect 83826 -90447 83904 -90442
rect 83478 -90930 83538 -90449
rect 83834 -90930 83894 -90447
rect 54845 -91316 86391 -90930
rect 54849 -91555 86391 -91316
rect 54849 -91941 86399 -91555
<< via3 >>
rect 68314 -70126 68390 -70086
rect 68314 -71268 68320 -70126
rect 68320 -71268 68382 -70126
rect 68382 -71268 68390 -70126
rect 68666 -70122 68742 -70086
rect 68666 -71266 68670 -70122
rect 68670 -71266 68732 -70122
rect 68732 -71266 68742 -70122
rect 68666 -71268 68742 -71266
rect 69020 -70116 69096 -70078
rect 69020 -71260 69026 -70116
rect 69026 -71260 69088 -70116
rect 69088 -71260 69096 -70116
rect 69376 -70120 69452 -70080
rect 69376 -71262 69378 -70120
rect 69378 -71262 69440 -70120
rect 69440 -71262 69452 -70120
rect 69728 -70118 69804 -70080
rect 69728 -71262 69732 -70118
rect 69732 -71262 69794 -70118
rect 69794 -71262 69804 -70118
rect 70090 -70122 70166 -70092
rect 70090 -71266 70094 -70122
rect 70094 -71266 70156 -70122
rect 70156 -71266 70166 -70122
rect 70090 -71274 70166 -71266
rect 70444 -70114 70520 -70078
rect 70444 -71258 70452 -70114
rect 70452 -71258 70514 -70114
rect 70514 -71258 70520 -70114
rect 70444 -71260 70520 -71258
rect 70792 -70110 70868 -70070
rect 70792 -71252 70804 -70110
rect 70804 -71252 70866 -70110
rect 70866 -71252 70868 -70110
rect 71150 -70114 71226 -70078
rect 71150 -71258 71158 -70114
rect 71158 -71258 71220 -70114
rect 71220 -71258 71226 -70114
rect 71150 -71260 71226 -71258
rect 71506 -70114 71582 -70080
rect 71506 -71258 71512 -70114
rect 71512 -71258 71574 -70114
rect 71574 -71258 71582 -70114
rect 71506 -71262 71582 -71258
rect 71868 -70114 71944 -70078
rect 71868 -71258 71874 -70114
rect 71874 -71258 71936 -70114
rect 71936 -71258 71944 -70114
rect 71868 -71260 71944 -71258
rect 72222 -70118 72298 -70078
rect 72222 -71260 72228 -70118
rect 72228 -71260 72290 -70118
rect 72290 -71260 72298 -70118
rect 72584 -70118 72660 -70074
rect 72584 -71256 72586 -70118
rect 72586 -71256 72648 -70118
rect 72648 -71256 72660 -70118
rect 72938 -70114 73014 -70076
rect 72938 -71258 72942 -70114
rect 72942 -71258 73004 -70114
rect 73004 -71258 73014 -70114
rect 73292 -70114 73368 -70078
rect 73292 -71258 73302 -70114
rect 73302 -71258 73364 -70114
rect 73364 -71258 73368 -70114
rect 73292 -71260 73368 -71258
rect 73642 -70118 73718 -70080
rect 73642 -71262 73652 -70118
rect 73652 -71262 73714 -70118
rect 73714 -71262 73718 -70118
rect 74004 -70114 74080 -70080
rect 74004 -71258 74008 -70114
rect 74008 -71258 74070 -70114
rect 74070 -71258 74080 -70114
rect 74004 -71262 74080 -71258
rect 74356 -70112 74432 -70074
rect 74356 -71256 74366 -70112
rect 74366 -71256 74428 -70112
rect 74428 -71256 74432 -70112
rect 74720 -70114 74796 -70084
rect 74720 -71258 74724 -70114
rect 74724 -71258 74786 -70114
rect 74786 -71258 74796 -70114
rect 74720 -71266 74796 -71258
rect 75070 -70114 75146 -70078
rect 75070 -71258 75074 -70114
rect 75074 -71258 75136 -70114
rect 75136 -71258 75146 -70114
rect 75070 -71260 75146 -71258
rect 75428 -70112 75504 -70078
rect 75428 -71256 75432 -70112
rect 75432 -71256 75494 -70112
rect 75494 -71256 75504 -70112
rect 75428 -71260 75504 -71256
rect 75782 -70112 75858 -70078
rect 75782 -71256 75788 -70112
rect 75788 -71256 75850 -70112
rect 75850 -71256 75858 -70112
rect 75782 -71260 75858 -71256
rect 76136 -70114 76212 -70078
rect 76136 -71258 76146 -70114
rect 76146 -71258 76208 -70114
rect 76208 -71258 76212 -70114
rect 76136 -71260 76212 -71258
rect 76492 -70112 76568 -70076
rect 76492 -71256 76496 -70112
rect 76496 -71256 76558 -70112
rect 76558 -71256 76568 -70112
rect 76492 -71258 76568 -71256
rect 76854 -70114 76930 -70088
rect 76854 -71258 76860 -70114
rect 76860 -71258 76922 -70114
rect 76922 -71258 76930 -70114
rect 76854 -71270 76930 -71258
rect 77198 -70118 77274 -70080
rect 77198 -71262 77212 -70118
rect 77212 -71262 77274 -70118
rect 77554 -70112 77630 -70080
rect 77554 -71256 77568 -70112
rect 77568 -71256 77630 -70112
rect 77554 -71262 77630 -71256
rect 77918 -70110 77994 -70074
rect 77918 -71254 77926 -70110
rect 77926 -71254 77988 -70110
rect 77988 -71254 77994 -70110
rect 77918 -71256 77994 -71254
rect 78272 -70112 78348 -70084
rect 78272 -71256 78282 -70112
rect 78282 -71256 78344 -70112
rect 78344 -71256 78348 -70112
rect 78272 -71266 78348 -71256
rect 78634 -70112 78710 -70080
rect 78634 -71256 78638 -70112
rect 78638 -71256 78700 -70112
rect 78700 -71256 78710 -70112
rect 78634 -71262 78710 -71256
rect 78992 -70114 79068 -70080
rect 78992 -71258 78996 -70114
rect 78996 -71258 79058 -70114
rect 79058 -71258 79068 -70114
rect 78992 -71262 79068 -71258
rect 79346 -70118 79422 -70084
rect 79346 -71262 79408 -70118
rect 79408 -71262 79422 -70118
rect 79346 -71266 79422 -71262
rect 79696 -70118 79772 -70078
rect 79696 -71260 79704 -70118
rect 79704 -71260 79766 -70118
rect 79766 -71260 79772 -70118
rect 80052 -70112 80128 -70084
rect 80052 -71256 80058 -70112
rect 80058 -71256 80120 -70112
rect 80120 -71256 80128 -70112
rect 80052 -71266 80128 -71256
rect 80412 -70118 80488 -70080
rect 80412 -71262 80474 -70118
rect 80474 -71262 80488 -70118
rect 80760 -70114 80836 -70080
rect 80760 -71258 80768 -70114
rect 80768 -71258 80830 -70114
rect 80830 -71258 80836 -70114
rect 80760 -71262 80836 -71258
rect 81114 -70118 81190 -70078
rect 81114 -71260 81126 -70118
rect 81126 -71260 81188 -70118
rect 81188 -71260 81190 -70118
rect 81478 -70114 81554 -70084
rect 81478 -71258 81480 -70114
rect 81480 -71258 81542 -70114
rect 81542 -71258 81554 -70114
rect 81478 -71266 81554 -71258
rect 81830 -70118 81906 -70080
rect 81830 -71262 81836 -70118
rect 81836 -71262 81898 -70118
rect 81898 -71262 81906 -70118
rect 82176 -70114 82252 -70080
rect 82176 -71258 82190 -70114
rect 82190 -71258 82252 -70114
rect 82176 -71262 82252 -71258
rect 82534 -70118 82610 -70086
rect 82534 -71262 82546 -70118
rect 82546 -71262 82608 -70118
rect 82608 -71262 82610 -70118
rect 82534 -71268 82610 -71262
rect 82894 -70114 82970 -70084
rect 82894 -71258 82906 -70114
rect 82906 -71258 82968 -70114
rect 82968 -71258 82970 -70114
rect 82894 -71266 82970 -71258
rect 83264 -70112 83340 -70070
rect 83264 -71252 83326 -70112
rect 83326 -71252 83340 -70112
rect 83616 -70118 83692 -70086
rect 83616 -71262 83620 -70118
rect 83620 -71262 83682 -70118
rect 83682 -71262 83692 -70118
rect 83616 -71268 83692 -71262
rect 83980 -70118 84056 -70086
rect 83980 -71262 84038 -70118
rect 84038 -71262 84056 -70118
rect 83980 -71268 84056 -71262
rect 68312 -71562 68376 -71542
rect 68312 -72676 68314 -71562
rect 68314 -72676 68376 -71562
rect 68662 -71540 68726 -71526
rect 68662 -72660 68664 -71540
rect 68664 -72660 68726 -71540
rect 69018 -71542 69082 -71526
rect 69018 -72652 69080 -71542
rect 69080 -72652 69082 -71542
rect 69018 -72660 69082 -72652
rect 69376 -71540 69440 -71526
rect 69376 -72660 69378 -71540
rect 69378 -72660 69440 -71540
rect 69724 -71548 69788 -71530
rect 69724 -72658 69786 -71548
rect 69786 -72658 69788 -71548
rect 69724 -72664 69788 -72658
rect 70088 -71536 70152 -71518
rect 70088 -72646 70148 -71536
rect 70148 -72646 70152 -71536
rect 70088 -72652 70152 -72646
rect 70450 -71542 70514 -71526
rect 70450 -72652 70512 -71542
rect 70512 -72652 70514 -71542
rect 70450 -72660 70514 -72652
rect 70790 -71546 70854 -71530
rect 70790 -72656 70852 -71546
rect 70852 -72656 70854 -71546
rect 70790 -72664 70854 -72656
rect 71148 -71554 71212 -71538
rect 71148 -72664 71210 -71554
rect 71210 -72664 71212 -71554
rect 71148 -72672 71212 -72664
rect 71504 -71546 71568 -71530
rect 71504 -72656 71566 -71546
rect 71566 -72656 71568 -71546
rect 71504 -72664 71568 -72656
rect 71858 -71542 71922 -71526
rect 71858 -72652 71920 -71542
rect 71920 -72652 71922 -71542
rect 71858 -72660 71922 -72652
rect 72218 -71546 72282 -71530
rect 72218 -72656 72278 -71546
rect 72278 -72656 72282 -71546
rect 72218 -72664 72282 -72656
rect 72572 -71544 72636 -71530
rect 72572 -72654 72632 -71544
rect 72632 -72654 72636 -71544
rect 72572 -72664 72636 -72654
rect 72944 -71542 73008 -71530
rect 72944 -72652 72946 -71542
rect 72946 -72652 73008 -71542
rect 72944 -72664 73008 -72652
rect 73286 -71558 73350 -71542
rect 73286 -72668 73348 -71558
rect 73348 -72668 73350 -71558
rect 73286 -72676 73350 -72668
rect 73642 -71550 73706 -71526
rect 73642 -72660 73704 -71550
rect 73704 -72660 73706 -71550
rect 73988 -71542 74052 -71518
rect 73988 -72652 74050 -71542
rect 74050 -72652 74052 -71542
rect 74352 -71560 74416 -71538
rect 74352 -72670 74414 -71560
rect 74414 -72670 74416 -71560
rect 74352 -72672 74416 -72670
rect 74714 -71556 74778 -71530
rect 74714 -72664 74776 -71556
rect 74776 -72664 74778 -71556
rect 75070 -71572 75134 -71550
rect 75070 -72682 75130 -71572
rect 75130 -72682 75134 -71572
rect 75070 -72684 75134 -72682
rect 75426 -71560 75490 -71538
rect 75426 -72670 75488 -71560
rect 75488 -72670 75490 -71560
rect 75426 -72672 75490 -72670
rect 75764 -71544 75828 -71518
rect 75764 -72652 75826 -71544
rect 75826 -72652 75828 -71544
rect 76128 -71542 76192 -71518
rect 76128 -72652 76130 -71542
rect 76130 -72652 76192 -71542
rect 76478 -71542 76542 -71518
rect 76478 -72652 76540 -71542
rect 76540 -72652 76542 -71542
rect 76854 -71546 76918 -71526
rect 76854 -72656 76916 -71546
rect 76916 -72656 76918 -71546
rect 76854 -72660 76918 -72656
rect 77196 -71550 77260 -71526
rect 77196 -72660 77258 -71550
rect 77258 -72660 77260 -71550
rect 77910 -71538 77974 -71514
rect 77548 -71562 77612 -71538
rect 77548 -72672 77610 -71562
rect 77610 -72672 77612 -71562
rect 77910 -72648 77970 -71538
rect 77970 -72648 77974 -71538
rect 78274 -71540 78338 -71518
rect 78274 -72650 78336 -71540
rect 78336 -72650 78338 -71540
rect 78274 -72652 78338 -72650
rect 78624 -71562 78688 -71538
rect 78624 -72672 78686 -71562
rect 78686 -72672 78688 -71562
rect 78988 -71562 79052 -71542
rect 78988 -72672 78990 -71562
rect 78990 -72672 79052 -71562
rect 78988 -72676 79052 -72672
rect 79338 -71542 79402 -71518
rect 79338 -72652 79400 -71542
rect 79400 -72652 79402 -71542
rect 79694 -71550 79758 -71526
rect 79694 -72660 79754 -71550
rect 79754 -72660 79758 -71550
rect 80046 -71556 80110 -71530
rect 80046 -72664 80048 -71556
rect 80048 -72664 80110 -71556
rect 80400 -71560 80464 -71538
rect 80400 -72670 80460 -71560
rect 80460 -72670 80464 -71560
rect 80400 -72672 80464 -72670
rect 80760 -71552 80824 -71526
rect 80760 -72660 80822 -71552
rect 80822 -72660 80824 -71552
rect 81122 -71562 81186 -71538
rect 81122 -72672 81182 -71562
rect 81182 -72672 81186 -71562
rect 81478 -71550 81542 -71530
rect 81478 -72660 81540 -71550
rect 81540 -72660 81542 -71550
rect 81478 -72664 81542 -72660
rect 81848 -71552 81912 -71530
rect 81848 -72662 81910 -71552
rect 81910 -72662 81912 -71552
rect 81848 -72664 81912 -72662
rect 82184 -71560 82248 -71538
rect 82184 -72670 82186 -71560
rect 82186 -72670 82248 -71560
rect 82184 -72672 82248 -72670
rect 82542 -71566 82606 -71542
rect 82542 -72676 82604 -71566
rect 82604 -72676 82606 -71566
rect 82906 -71574 82970 -71550
rect 82906 -72684 82910 -71574
rect 82910 -72684 82970 -71574
rect 83256 -71552 83320 -71530
rect 83256 -72662 83258 -71552
rect 83258 -72662 83320 -71552
rect 83256 -72664 83320 -72662
rect 83612 -71574 83676 -71550
rect 83612 -72684 83674 -71574
rect 83674 -72684 83676 -71574
rect 83962 -71550 84026 -71530
rect 83962 -72660 84024 -71550
rect 84024 -72660 84026 -71550
rect 83962 -72664 84026 -72660
rect 56466 -74540 56488 -73428
rect 56488 -74540 56544 -73428
rect 56544 -74540 56560 -73428
rect 56854 -74534 56908 -73428
rect 56908 -74534 56948 -73428
rect 56466 -74542 56560 -74540
rect 56854 -74542 56948 -74534
rect 57186 -74542 57196 -73428
rect 57196 -74542 57252 -73428
rect 57252 -74542 57280 -73428
rect 57542 -74526 57556 -73412
rect 57556 -74526 57612 -73412
rect 57612 -74526 57636 -73412
rect 57890 -74536 57916 -73422
rect 57916 -74536 57972 -73422
rect 57972 -74536 57984 -73422
rect 58256 -74526 58274 -73412
rect 58274 -74526 58330 -73412
rect 58330 -74526 58350 -73412
rect 58616 -74526 58628 -73412
rect 58628 -74526 58684 -73412
rect 58684 -74526 58710 -73412
rect 58970 -74542 58980 -73428
rect 58980 -74542 59036 -73428
rect 59036 -74542 59064 -73428
rect 59330 -74538 59342 -73428
rect 59342 -74538 59398 -73428
rect 59398 -74538 59424 -73428
rect 59672 -74536 59694 -73422
rect 59694 -74536 59750 -73422
rect 59750 -74536 59766 -73422
rect 59330 -74542 59424 -74538
rect 56468 -75988 56472 -74874
rect 56472 -75988 56528 -74874
rect 56528 -75988 56562 -74874
rect 56828 -75988 56836 -74874
rect 56836 -75988 56892 -74874
rect 56892 -75988 56922 -74874
rect 57178 -75998 57180 -74884
rect 57180 -75998 57236 -74884
rect 57236 -75998 57272 -74884
rect 57532 -75988 57540 -74874
rect 57540 -75988 57596 -74874
rect 57596 -75988 57626 -74874
rect 57896 -75998 57900 -74884
rect 57900 -75998 57956 -74884
rect 57956 -75998 57990 -74884
rect 58246 -75988 58258 -74874
rect 58258 -75988 58314 -74874
rect 58314 -75988 58340 -74874
rect 58600 -75982 58612 -74868
rect 58612 -75982 58668 -74868
rect 58668 -75982 58694 -74868
rect 58960 -75988 58964 -74874
rect 58964 -75988 59020 -74874
rect 59020 -75988 59054 -74874
rect 59320 -75982 59326 -74868
rect 59326 -75982 59382 -74868
rect 59382 -75982 59414 -74868
rect 59668 -75998 59678 -74884
rect 59678 -75998 59734 -74884
rect 59734 -75998 59762 -74884
rect 56456 -78390 56478 -77284
rect 56478 -78390 56534 -77284
rect 56534 -78390 56550 -77284
rect 56456 -78398 56550 -78390
rect 56816 -78384 56842 -77284
rect 56842 -78384 56898 -77284
rect 56898 -78384 56910 -77284
rect 56816 -78398 56910 -78384
rect 57166 -78396 57186 -77294
rect 57186 -78396 57242 -77294
rect 57242 -78396 57260 -77294
rect 57166 -78408 57260 -78396
rect 57520 -78390 57546 -77284
rect 57546 -78390 57602 -77284
rect 57602 -78390 57614 -77284
rect 57520 -78398 57614 -78390
rect 57884 -78396 57906 -77294
rect 57906 -78396 57962 -77294
rect 57962 -78396 57978 -77294
rect 57884 -78408 57978 -78396
rect 58234 -78398 58264 -77284
rect 58264 -78398 58320 -77284
rect 58320 -78398 58328 -77284
rect 58588 -78388 58618 -77278
rect 58618 -78388 58674 -77278
rect 58674 -78388 58682 -77278
rect 58588 -78392 58682 -78388
rect 58948 -78392 58970 -77284
rect 58970 -78392 59026 -77284
rect 59026 -78392 59042 -77284
rect 59308 -78388 59332 -77278
rect 59332 -78388 59388 -77278
rect 59388 -78388 59402 -77278
rect 59308 -78392 59402 -78388
rect 59656 -78392 59684 -77294
rect 59684 -78392 59740 -77294
rect 59740 -78392 59750 -77294
rect 58948 -78398 59042 -78392
rect 59656 -78408 59750 -78392
rect 56440 -79834 56462 -78720
rect 56462 -79834 56518 -78720
rect 56518 -79834 56534 -78720
rect 56800 -79834 56826 -78720
rect 56826 -79834 56882 -78720
rect 56882 -79834 56894 -78720
rect 57150 -79844 57170 -78730
rect 57170 -79844 57226 -78730
rect 57226 -79844 57244 -78730
rect 57504 -79834 57530 -78720
rect 57530 -79834 57586 -78720
rect 57586 -79834 57598 -78720
rect 58218 -78722 58312 -78720
rect 57868 -79844 57890 -78730
rect 57890 -79844 57946 -78730
rect 57946 -79844 57962 -78730
rect 58218 -79834 58248 -78722
rect 58248 -79834 58304 -78722
rect 58304 -79834 58312 -78722
rect 58572 -79828 58602 -78714
rect 58602 -79828 58658 -78714
rect 58658 -79828 58666 -78714
rect 58932 -79834 58954 -78720
rect 58954 -79834 59010 -78720
rect 59010 -79834 59026 -78720
rect 59292 -79828 59316 -78714
rect 59316 -79828 59372 -78714
rect 59372 -79828 59386 -78714
rect 59640 -79844 59668 -78730
rect 59668 -79844 59724 -78730
rect 59724 -79844 59734 -78730
rect 61102 -82360 61118 -81246
rect 61118 -82360 61174 -81246
rect 61174 -82360 61196 -81246
rect 61462 -82344 61476 -81230
rect 61476 -82344 61532 -81230
rect 61532 -82344 61556 -81230
rect 61810 -82344 61826 -81230
rect 61826 -82344 61882 -81230
rect 61882 -82344 61904 -81230
rect 62170 -82344 62188 -81230
rect 62188 -82344 62244 -81230
rect 62244 -82344 62264 -81230
rect 62530 -82350 62544 -81236
rect 62544 -82350 62600 -81236
rect 62600 -82350 62624 -81236
rect 62884 -82350 62894 -81236
rect 62894 -82350 62950 -81236
rect 62950 -82350 62978 -81236
rect 63234 -82350 63254 -81236
rect 63254 -82350 63310 -81236
rect 63310 -82350 63328 -81236
rect 63594 -82360 63614 -81246
rect 63614 -82360 63670 -81246
rect 63670 -82360 63688 -81246
rect 63952 -82344 63966 -81230
rect 63966 -82344 64022 -81230
rect 64022 -82344 64046 -81230
rect 64296 -82344 64320 -81230
rect 64320 -82344 64376 -81230
rect 64376 -82344 64390 -81230
rect 61444 -82682 61538 -82676
rect 61086 -83816 61102 -82702
rect 61102 -83816 61158 -82702
rect 61158 -83816 61180 -82702
rect 61444 -83790 61460 -82682
rect 61460 -83790 61516 -82682
rect 61516 -83790 61538 -82682
rect 61788 -82688 61882 -82676
rect 61788 -83790 61810 -82688
rect 61810 -83790 61866 -82688
rect 61866 -83790 61882 -82688
rect 62164 -82692 62258 -82676
rect 62164 -83790 62172 -82692
rect 62172 -83790 62228 -82692
rect 62228 -83790 62258 -82692
rect 62514 -82688 62608 -82676
rect 62514 -83790 62528 -82688
rect 62528 -83790 62584 -82688
rect 62584 -83790 62608 -82688
rect 62856 -82692 62950 -82686
rect 63576 -82692 63670 -82670
rect 62856 -83800 62878 -82692
rect 62878 -83800 62934 -82692
rect 62934 -83800 62950 -82692
rect 63216 -83806 63238 -82692
rect 63238 -83806 63294 -82692
rect 63294 -83806 63310 -82692
rect 63576 -83784 63598 -82692
rect 63598 -83784 63654 -82692
rect 63654 -83784 63670 -82692
rect 63920 -83800 63950 -82686
rect 63950 -83800 64006 -82686
rect 64006 -83800 64014 -82686
rect 64286 -83806 64304 -82692
rect 64304 -83806 64360 -82692
rect 64360 -83806 64380 -82692
rect 61778 -85046 61872 -85036
rect 61068 -86182 61090 -85068
rect 61090 -86182 61146 -85068
rect 61146 -86182 61162 -85068
rect 61418 -86160 61448 -85046
rect 61448 -86160 61504 -85046
rect 61504 -86160 61512 -85046
rect 61778 -86150 61798 -85046
rect 61798 -86150 61854 -85046
rect 61854 -86150 61872 -85046
rect 62154 -85050 62248 -85036
rect 62154 -86150 62160 -85050
rect 62160 -86150 62216 -85050
rect 62216 -86150 62248 -85050
rect 62492 -85046 62586 -85036
rect 64270 -85044 64364 -85024
rect 62492 -86150 62516 -85046
rect 62516 -86150 62572 -85046
rect 62572 -86150 62586 -85046
rect 62840 -86178 62866 -85064
rect 62866 -86178 62922 -85064
rect 62922 -86178 62934 -85064
rect 63206 -86178 63226 -85064
rect 63226 -86178 63282 -85064
rect 63282 -86178 63300 -85064
rect 63566 -86166 63586 -85052
rect 63586 -86166 63642 -85052
rect 63642 -86166 63660 -85052
rect 63926 -86166 63938 -85052
rect 63938 -86166 63994 -85052
rect 63994 -86166 64020 -85052
rect 64270 -86138 64292 -85044
rect 64292 -86138 64348 -85044
rect 64348 -86138 64364 -85044
rect 61058 -86508 61152 -86480
rect 61058 -87594 61074 -86508
rect 61074 -87594 61130 -86508
rect 61130 -87594 61152 -86508
rect 61418 -86502 61512 -86498
rect 61418 -87612 61432 -86502
rect 61432 -87612 61488 -86502
rect 61488 -87612 61512 -86502
rect 62132 -86512 62226 -86498
rect 61772 -87632 61782 -86518
rect 61782 -87632 61838 -86518
rect 61838 -87632 61866 -86518
rect 62132 -87612 62144 -86512
rect 62144 -87612 62200 -86512
rect 62200 -87612 62226 -86512
rect 62492 -86508 62586 -86492
rect 62492 -87606 62500 -86508
rect 62500 -87606 62556 -86508
rect 62556 -87606 62586 -86508
rect 63200 -86510 63294 -86508
rect 62840 -87632 62850 -86518
rect 62850 -87632 62906 -86518
rect 62906 -87632 62934 -86518
rect 63200 -87622 63210 -86510
rect 63210 -87622 63266 -86510
rect 63266 -87622 63294 -86510
rect 63560 -86512 63654 -86498
rect 63560 -87612 63570 -86512
rect 63570 -87612 63626 -86512
rect 63626 -87612 63654 -86512
rect 63910 -87622 63922 -86508
rect 63922 -87622 63978 -86508
rect 63978 -87622 64004 -86508
rect 64270 -87622 64276 -86508
rect 64276 -87622 64332 -86508
rect 64332 -87622 64364 -86508
rect 68436 -89014 68440 -87882
rect 68440 -89014 68498 -87882
rect 68498 -89014 68504 -87882
rect 68798 -89022 68802 -87890
rect 68802 -89022 68860 -87890
rect 68860 -89022 68866 -87890
rect 69148 -89022 69160 -87890
rect 69160 -89022 69216 -87890
rect 56534 -90468 56542 -89346
rect 56542 -90468 56602 -89346
rect 56602 -90468 56610 -89346
rect 56894 -90464 56900 -89342
rect 56900 -90464 56960 -89342
rect 56960 -90464 56970 -89342
rect 57250 -90474 57254 -89352
rect 57254 -90474 57314 -89352
rect 57314 -90474 57326 -89352
rect 57600 -90474 57608 -89352
rect 57608 -90474 57668 -89352
rect 57668 -90474 57676 -89352
rect 57956 -90472 57964 -89350
rect 57964 -90472 58024 -89350
rect 58024 -90472 58032 -89350
rect 58312 -90470 58322 -89348
rect 58322 -90470 58382 -89348
rect 58382 -90470 58388 -89348
rect 58674 -90460 58682 -89338
rect 58682 -90460 58742 -89338
rect 58742 -90460 58750 -89338
rect 59024 -90472 59028 -89350
rect 59028 -90472 59088 -89350
rect 59088 -90472 59100 -89350
rect 59386 -90462 59388 -89340
rect 59388 -90462 59448 -89340
rect 59448 -90462 59462 -89340
rect 59736 -90456 59746 -89334
rect 59746 -90456 59806 -89334
rect 59806 -90456 59812 -89334
rect 60964 -90464 60974 -89342
rect 60974 -90464 61034 -89342
rect 61034 -90464 61040 -89342
rect 61318 -90474 61322 -89352
rect 61322 -90474 61382 -89352
rect 61382 -90474 61394 -89352
rect 61676 -90460 61680 -89338
rect 61680 -90460 61740 -89338
rect 61740 -90460 61752 -89338
rect 62036 -90470 62042 -89348
rect 62042 -90470 62102 -89348
rect 62102 -90470 62112 -89348
rect 62392 -90476 62396 -89354
rect 62396 -90476 62456 -89354
rect 62456 -90476 62468 -89354
rect 62742 -90474 62752 -89352
rect 62752 -90474 62812 -89352
rect 62812 -90474 62818 -89352
rect 63104 -90468 63106 -89346
rect 63106 -90468 63166 -89346
rect 63166 -90468 63180 -89346
rect 63458 -90482 63466 -89360
rect 63466 -90482 63526 -89360
rect 63526 -90482 63534 -89360
rect 63816 -90468 63826 -89346
rect 63826 -90468 63886 -89346
rect 63886 -90468 63892 -89346
rect 64176 -90474 64182 -89352
rect 64182 -90474 64242 -89352
rect 64242 -90474 64252 -89352
rect 68440 -90440 68444 -89308
rect 68444 -90440 68502 -89308
rect 68502 -90440 68508 -89308
rect 69506 -89024 69512 -87892
rect 69512 -89024 69570 -87892
rect 69570 -89024 69574 -87892
rect 69860 -89020 69866 -87888
rect 69866 -89020 69924 -87888
rect 69924 -89020 69928 -87888
rect 68796 -90440 68800 -89308
rect 68800 -90440 68858 -89308
rect 68858 -90440 68864 -89308
rect 70212 -89026 70222 -87894
rect 70222 -89026 70280 -87894
rect 70574 -89022 70582 -87890
rect 70582 -89022 70640 -87890
rect 70640 -89022 70642 -87890
rect 69150 -90440 69156 -89308
rect 69156 -90440 69214 -89308
rect 69214 -90440 69218 -89308
rect 69500 -90442 69508 -89310
rect 69508 -90442 69566 -89310
rect 69566 -90442 69568 -89310
rect 69856 -90448 69864 -89316
rect 69864 -90448 69922 -89316
rect 69922 -90448 69924 -89316
rect 70928 -89026 70936 -87894
rect 70936 -89026 70994 -87894
rect 70994 -89026 70996 -87894
rect 71286 -89030 71292 -87898
rect 71292 -89030 71350 -87898
rect 71350 -89030 71354 -87898
rect 71644 -89026 71646 -87894
rect 71646 -89026 71704 -87894
rect 71704 -89026 71712 -87894
rect 74332 -89012 74336 -87880
rect 74336 -89012 74394 -87880
rect 74394 -89012 74400 -87880
rect 74694 -89020 74698 -87888
rect 74698 -89020 74756 -87888
rect 74756 -89020 74762 -87888
rect 70220 -90444 70226 -89316
rect 70226 -90444 70284 -89316
rect 70284 -90444 70288 -89316
rect 70220 -90448 70288 -90444
rect 70570 -90446 70578 -89314
rect 70578 -90446 70636 -89314
rect 70636 -90446 70638 -89314
rect 70926 -90444 70934 -89312
rect 70934 -90444 70992 -89312
rect 70992 -90444 70994 -89312
rect 71286 -90448 71294 -89316
rect 71294 -90448 71352 -89316
rect 71352 -90448 71354 -89316
rect 71634 -90446 71646 -89316
rect 71646 -90446 71702 -89316
rect 71634 -90448 71702 -90446
rect 75044 -89020 75056 -87888
rect 75056 -89020 75112 -87888
rect 74336 -90438 74340 -89306
rect 74340 -90438 74398 -89306
rect 74398 -90438 74404 -89306
rect 75402 -89022 75408 -87890
rect 75408 -89022 75466 -87890
rect 75466 -89022 75470 -87890
rect 75756 -89018 75762 -87886
rect 75762 -89018 75820 -87886
rect 75820 -89018 75824 -87886
rect 74692 -90438 74696 -89306
rect 74696 -90438 74754 -89306
rect 74754 -90438 74760 -89306
rect 75046 -90438 75052 -89306
rect 75052 -90438 75110 -89306
rect 75110 -90438 75114 -89306
rect 76108 -89024 76118 -87892
rect 76118 -89024 76176 -87892
rect 76470 -89020 76478 -87888
rect 76478 -89020 76536 -87888
rect 76536 -89020 76538 -87888
rect 75396 -90440 75404 -89308
rect 75404 -90440 75462 -89308
rect 75462 -90440 75464 -89308
rect 75752 -90446 75760 -89314
rect 75760 -90446 75818 -89314
rect 75818 -90446 75820 -89314
rect 76824 -89024 76832 -87892
rect 76832 -89024 76890 -87892
rect 76890 -89024 76892 -87892
rect 77182 -89028 77188 -87896
rect 77188 -89028 77246 -87896
rect 77246 -89028 77250 -87896
rect 77540 -89024 77542 -87892
rect 77542 -89024 77600 -87892
rect 77600 -89024 77608 -87892
rect 80446 -89006 80450 -87874
rect 80450 -89006 80508 -87874
rect 80508 -89006 80514 -87874
rect 80808 -89014 80812 -87882
rect 80812 -89014 80870 -87882
rect 80870 -89014 80876 -87882
rect 76116 -90442 76122 -89314
rect 76122 -90442 76180 -89314
rect 76180 -90442 76184 -89314
rect 76116 -90446 76184 -90442
rect 76466 -90444 76474 -89312
rect 76474 -90444 76532 -89312
rect 76532 -90444 76534 -89312
rect 76822 -90442 76830 -89310
rect 76830 -90442 76888 -89310
rect 76888 -90442 76890 -89310
rect 77182 -90446 77190 -89314
rect 77190 -90446 77248 -89314
rect 77248 -90446 77250 -89314
rect 77530 -90444 77542 -89314
rect 77542 -90444 77598 -89314
rect 77530 -90446 77598 -90444
rect 81158 -89014 81170 -87882
rect 81170 -89014 81226 -87882
rect 80450 -90432 80454 -89300
rect 80454 -90432 80512 -89300
rect 80512 -90432 80518 -89300
rect 81516 -89016 81522 -87884
rect 81522 -89016 81580 -87884
rect 81580 -89016 81584 -87884
rect 81870 -89012 81876 -87880
rect 81876 -89012 81934 -87880
rect 81934 -89012 81938 -87880
rect 80806 -90432 80810 -89300
rect 80810 -90432 80868 -89300
rect 80868 -90432 80874 -89300
rect 82222 -89018 82232 -87886
rect 82232 -89018 82290 -87886
rect 82584 -89014 82592 -87882
rect 82592 -89014 82650 -87882
rect 82650 -89014 82652 -87882
rect 81160 -90432 81166 -89300
rect 81166 -90432 81224 -89300
rect 81224 -90432 81228 -89300
rect 81510 -90434 81518 -89302
rect 81518 -90434 81576 -89302
rect 81576 -90434 81578 -89302
rect 81866 -90440 81874 -89308
rect 81874 -90440 81932 -89308
rect 81932 -90440 81934 -89308
rect 82938 -89018 82946 -87886
rect 82946 -89018 83004 -87886
rect 83004 -89018 83006 -87886
rect 83296 -89022 83302 -87890
rect 83302 -89022 83360 -87890
rect 83360 -89022 83364 -87890
rect 83654 -89018 83656 -87886
rect 83656 -89018 83714 -87886
rect 83714 -89018 83722 -87886
rect 82230 -90436 82236 -89308
rect 82236 -90436 82294 -89308
rect 82294 -90436 82298 -89308
rect 82230 -90440 82298 -90436
rect 82580 -90438 82588 -89306
rect 82588 -90438 82646 -89306
rect 82646 -90438 82648 -89306
rect 82936 -90436 82944 -89304
rect 82944 -90436 83002 -89304
rect 83002 -90436 83004 -89304
rect 83296 -90440 83304 -89308
rect 83304 -90440 83362 -89308
rect 83362 -90440 83364 -89308
rect 83644 -90438 83656 -89308
rect 83656 -90438 83712 -89308
rect 83644 -90440 83712 -90438
<< metal4 >>
rect 56240 -73412 60060 -73348
rect 56240 -73428 57542 -73412
rect 56240 -74542 56466 -73428
rect 56560 -74542 56854 -73428
rect 56948 -74542 57186 -73428
rect 57280 -74526 57542 -73428
rect 57636 -73422 58256 -73412
rect 57636 -74526 57890 -73422
rect 57280 -74536 57890 -74526
rect 57984 -74526 58256 -73422
rect 58350 -74526 58616 -73412
rect 58710 -73422 60060 -73412
rect 58710 -73428 59672 -73422
rect 58710 -74526 58970 -73428
rect 57984 -74536 58970 -74526
rect 57280 -74542 58970 -74536
rect 59064 -74542 59330 -73428
rect 59424 -74536 59672 -73428
rect 59766 -74536 60060 -73422
rect 59424 -74542 60060 -74536
rect 56240 -74868 60060 -74542
rect 56240 -74874 58600 -74868
rect 56240 -75988 56468 -74874
rect 56562 -75988 56828 -74874
rect 56922 -74884 57532 -74874
rect 56922 -75988 57178 -74884
rect 56240 -75998 57178 -75988
rect 57272 -75988 57532 -74884
rect 57626 -74884 58246 -74874
rect 57626 -75988 57896 -74884
rect 57272 -75998 57896 -75988
rect 57990 -75988 58246 -74884
rect 58340 -75982 58600 -74874
rect 58694 -74874 59320 -74868
rect 58694 -75982 58960 -74874
rect 58340 -75988 58960 -75982
rect 59054 -75982 59320 -74874
rect 59414 -74884 60060 -74868
rect 59414 -75982 59668 -74884
rect 59054 -75988 59668 -75982
rect 57990 -75998 59668 -75988
rect 59762 -75998 60060 -74884
rect 56240 -77278 60060 -75998
rect 56240 -77284 58588 -77278
rect 56240 -78398 56456 -77284
rect 56550 -78398 56816 -77284
rect 56910 -77294 57520 -77284
rect 56910 -78398 57166 -77294
rect 56240 -78408 57166 -78398
rect 57260 -78398 57520 -77294
rect 57614 -77294 58234 -77284
rect 57614 -78398 57884 -77294
rect 57260 -78408 57884 -78398
rect 57978 -78398 58234 -77294
rect 58328 -78392 58588 -77284
rect 58682 -77284 59308 -77278
rect 58682 -78392 58948 -77284
rect 58328 -78398 58948 -78392
rect 59042 -78392 59308 -77284
rect 59402 -77294 60060 -77278
rect 59402 -78392 59656 -77294
rect 59042 -78398 59656 -78392
rect 57978 -78408 59656 -78398
rect 59750 -78408 60060 -77294
rect 56240 -78714 60060 -78408
rect 56240 -78720 58572 -78714
rect 56240 -79834 56440 -78720
rect 56534 -79834 56800 -78720
rect 56894 -78730 57504 -78720
rect 56894 -79834 57150 -78730
rect 56240 -79844 57150 -79834
rect 57244 -79834 57504 -78730
rect 57598 -78730 58218 -78720
rect 57598 -79834 57868 -78730
rect 57244 -79844 57868 -79834
rect 57962 -79834 58218 -78730
rect 58312 -79828 58572 -78720
rect 58666 -78720 59292 -78714
rect 58666 -79828 58932 -78720
rect 58312 -79834 58932 -79828
rect 59026 -79828 59292 -78720
rect 59386 -78730 60060 -78714
rect 59386 -79828 59640 -78730
rect 59026 -79834 59640 -79828
rect 57962 -79844 59640 -79834
rect 59734 -79844 60060 -78730
rect 56240 -89334 60060 -79844
rect 60748 -81230 64462 -81046
rect 60748 -81246 61462 -81230
rect 60748 -82360 61102 -81246
rect 61196 -82344 61462 -81246
rect 61556 -82344 61810 -81230
rect 61904 -82344 62170 -81230
rect 62264 -81236 63952 -81230
rect 62264 -82344 62530 -81236
rect 61196 -82350 62530 -82344
rect 62624 -82350 62884 -81236
rect 62978 -82350 63234 -81236
rect 63328 -81246 63952 -81236
rect 63328 -82350 63594 -81246
rect 61196 -82360 63594 -82350
rect 63688 -82344 63952 -81246
rect 64046 -82344 64296 -81230
rect 64390 -82344 64462 -81230
rect 63688 -82360 64462 -82344
rect 60748 -82670 64462 -82360
rect 60748 -82676 63576 -82670
rect 60748 -82702 61444 -82676
rect 60748 -83816 61086 -82702
rect 61180 -83790 61444 -82702
rect 61538 -83790 61788 -82676
rect 61882 -83790 62164 -82676
rect 62258 -83790 62514 -82676
rect 62608 -82686 63576 -82676
rect 62608 -83790 62856 -82686
rect 61180 -83800 62856 -83790
rect 62950 -82692 63576 -82686
rect 62950 -83800 63216 -82692
rect 61180 -83806 63216 -83800
rect 63310 -83784 63576 -82692
rect 63670 -82686 64462 -82670
rect 63670 -83784 63920 -82686
rect 63310 -83800 63920 -83784
rect 64014 -82692 64462 -82686
rect 64014 -83800 64286 -82692
rect 63310 -83806 64286 -83800
rect 64380 -83806 64462 -82692
rect 61180 -83816 64462 -83806
rect 60748 -83986 64462 -83816
rect 60712 -84928 64462 -83986
rect 60748 -85024 64462 -84928
rect 60748 -85036 64270 -85024
rect 60748 -85046 61778 -85036
rect 60748 -85068 61418 -85046
rect 60748 -86182 61068 -85068
rect 61162 -86160 61418 -85068
rect 61512 -86150 61778 -85046
rect 61872 -86150 62154 -85036
rect 62248 -86150 62492 -85036
rect 62586 -85052 64270 -85036
rect 62586 -85064 63566 -85052
rect 62586 -86150 62840 -85064
rect 61512 -86160 62840 -86150
rect 61162 -86178 62840 -86160
rect 62934 -86178 63206 -85064
rect 63300 -86166 63566 -85064
rect 63660 -86166 63926 -85052
rect 64020 -86138 64270 -85052
rect 64364 -86138 64462 -85024
rect 64020 -86166 64462 -86138
rect 63300 -86178 64462 -86166
rect 61162 -86182 64462 -86178
rect 60748 -86480 64462 -86182
rect 60748 -87594 61058 -86480
rect 61152 -86492 64462 -86480
rect 61152 -86498 62492 -86492
rect 61152 -87594 61418 -86498
rect 60748 -87612 61418 -87594
rect 61512 -86518 62132 -86498
rect 61512 -87612 61772 -86518
rect 60748 -87632 61772 -87612
rect 61866 -87612 62132 -86518
rect 62226 -87606 62492 -86498
rect 62586 -86498 64462 -86492
rect 62586 -86508 63560 -86498
rect 62586 -86518 63200 -86508
rect 62586 -87606 62840 -86518
rect 62226 -87612 62840 -87606
rect 61866 -87632 62840 -87612
rect 62934 -87622 63200 -86518
rect 63294 -87612 63560 -86508
rect 63654 -86508 64462 -86498
rect 63654 -87612 63910 -86508
rect 63294 -87622 63910 -87612
rect 64004 -87622 64270 -86508
rect 64364 -87622 64462 -86508
rect 65956 -87374 66516 -69290
rect 70791 -70070 70869 -70069
rect 68310 -70085 68370 -70074
rect 69019 -70078 69097 -70077
rect 68668 -70085 68728 -70080
rect 68310 -70086 68391 -70085
rect 68310 -71268 68314 -70086
rect 68390 -71268 68391 -70086
rect 68310 -71269 68391 -71268
rect 68665 -70086 68743 -70085
rect 68665 -71268 68666 -70086
rect 68742 -71268 68743 -70086
rect 69019 -71260 69020 -70078
rect 69096 -71260 69097 -70078
rect 69734 -70079 69794 -70074
rect 70446 -70077 70506 -70074
rect 70443 -70078 70521 -70077
rect 69019 -71261 69097 -71260
rect 69375 -70080 69453 -70079
rect 68665 -71269 68743 -71268
rect 68310 -71541 68370 -71269
rect 68668 -71525 68728 -71269
rect 69020 -71525 69080 -71261
rect 69375 -71262 69376 -70080
rect 69452 -71262 69453 -70080
rect 69375 -71263 69453 -71262
rect 69727 -70080 69805 -70079
rect 69727 -71262 69728 -70080
rect 69804 -71262 69805 -70080
rect 69727 -71263 69805 -71262
rect 70088 -70091 70148 -70078
rect 70088 -70092 70167 -70091
rect 69376 -71525 69436 -71263
rect 68661 -71526 68728 -71525
rect 68310 -71542 68377 -71541
rect 68310 -72676 68312 -71542
rect 68376 -72676 68377 -71542
rect 68661 -72660 68662 -71526
rect 68726 -72660 68728 -71526
rect 68661 -72661 68728 -72660
rect 69017 -71526 69083 -71525
rect 69017 -72660 69018 -71526
rect 69082 -72660 69083 -71526
rect 69017 -72661 69083 -72660
rect 69375 -71526 69441 -71525
rect 69375 -72660 69376 -71526
rect 69440 -72660 69441 -71526
rect 69734 -71529 69794 -71263
rect 70088 -71274 70090 -70092
rect 70166 -71274 70167 -70092
rect 70443 -71260 70444 -70078
rect 70520 -71260 70521 -70078
rect 70791 -71252 70792 -70070
rect 70868 -71252 70869 -70070
rect 83263 -70070 83341 -70069
rect 72583 -70074 72661 -70073
rect 71156 -70077 71216 -70074
rect 70791 -71253 70869 -71252
rect 71149 -70078 71227 -70077
rect 70443 -71261 70521 -71260
rect 70088 -71275 70167 -71274
rect 70088 -71517 70148 -71275
rect 69375 -72661 69441 -72660
rect 69723 -71530 69794 -71529
rect 68310 -72677 68377 -72676
rect 68310 -73704 68370 -72677
rect 68668 -73704 68728 -72661
rect 69020 -73704 69080 -72661
rect 69376 -73704 69436 -72661
rect 69723 -72664 69724 -71530
rect 69788 -72664 69794 -71530
rect 70087 -71518 70153 -71517
rect 70087 -72652 70088 -71518
rect 70152 -72652 70153 -71518
rect 70087 -72653 70153 -72652
rect 70446 -71525 70506 -71261
rect 70446 -71526 70515 -71525
rect 69723 -72665 69794 -72664
rect 69734 -73704 69794 -72665
rect 70088 -73704 70148 -72653
rect 70446 -72660 70450 -71526
rect 70514 -72660 70515 -71526
rect 70800 -71529 70860 -71253
rect 71149 -71260 71150 -70078
rect 71226 -71260 71227 -70078
rect 71867 -70078 71945 -70077
rect 71149 -71261 71227 -71260
rect 71505 -70080 71583 -70079
rect 70446 -72661 70515 -72660
rect 70789 -71530 70860 -71529
rect 70446 -73704 70506 -72661
rect 70789 -72664 70790 -71530
rect 70854 -72664 70860 -71530
rect 71156 -71537 71216 -71261
rect 71505 -71262 71506 -70080
rect 71582 -71262 71583 -70080
rect 71867 -71260 71868 -70078
rect 71944 -71260 71945 -70078
rect 71867 -71261 71945 -71260
rect 72221 -70078 72299 -70077
rect 72583 -70078 72584 -70074
rect 72221 -71260 72222 -70078
rect 72298 -71260 72299 -70078
rect 72221 -71261 72299 -71260
rect 72580 -71256 72584 -70078
rect 72660 -71256 72661 -70074
rect 74355 -70074 74433 -70073
rect 77917 -70074 77995 -70073
rect 72937 -70076 73015 -70075
rect 72937 -70080 72938 -70076
rect 72580 -71257 72661 -71256
rect 71505 -71263 71583 -71262
rect 71512 -71529 71572 -71263
rect 71868 -71525 71928 -71261
rect 70789 -72665 70860 -72664
rect 70800 -73704 70860 -72665
rect 71147 -71538 71216 -71537
rect 71147 -72672 71148 -71538
rect 71212 -72672 71216 -71538
rect 71503 -71530 71572 -71529
rect 71503 -72664 71504 -71530
rect 71568 -72664 71572 -71530
rect 71857 -71526 71928 -71525
rect 71857 -72660 71858 -71526
rect 71922 -72660 71928 -71526
rect 72224 -71529 72284 -71261
rect 72580 -71529 72640 -71257
rect 71857 -72661 71928 -72660
rect 71503 -72665 71572 -72664
rect 71147 -72673 71216 -72672
rect 71156 -73704 71216 -72673
rect 71512 -73704 71572 -72665
rect 71868 -73704 71928 -72661
rect 72217 -71530 72284 -71529
rect 72217 -72664 72218 -71530
rect 72282 -72664 72284 -71530
rect 72217 -72665 72284 -72664
rect 72571 -71530 72640 -71529
rect 72571 -72664 72572 -71530
rect 72636 -72664 72640 -71530
rect 72571 -72665 72640 -72664
rect 72224 -73704 72284 -72665
rect 72580 -73704 72640 -72665
rect 72936 -71258 72938 -70080
rect 73014 -71258 73015 -70076
rect 72936 -71259 73015 -71258
rect 73291 -70078 73369 -70077
rect 72936 -71529 72996 -71259
rect 73291 -71260 73292 -70078
rect 73368 -71260 73369 -70078
rect 73650 -70079 73710 -70078
rect 73291 -71261 73369 -71260
rect 73641 -70080 73719 -70079
rect 72936 -71530 73009 -71529
rect 72936 -72664 72944 -71530
rect 73008 -72664 73009 -71530
rect 73294 -71541 73354 -71261
rect 73641 -71262 73642 -70080
rect 73718 -71262 73719 -70080
rect 73641 -71263 73719 -71262
rect 74003 -70080 74081 -70079
rect 74003 -71262 74004 -70080
rect 74080 -71262 74081 -70080
rect 74355 -71256 74356 -70074
rect 74432 -71256 74433 -70074
rect 76491 -70076 76569 -70075
rect 75069 -70078 75147 -70077
rect 74355 -71257 74433 -71256
rect 74716 -70083 74776 -70078
rect 74716 -70084 74797 -70083
rect 74003 -71263 74081 -71262
rect 73650 -71525 73710 -71263
rect 74004 -71517 74064 -71263
rect 72936 -72665 73009 -72664
rect 73285 -71542 73354 -71541
rect 72936 -73704 72996 -72665
rect 73285 -72676 73286 -71542
rect 73350 -72676 73354 -71542
rect 73641 -71526 73710 -71525
rect 73641 -72660 73642 -71526
rect 73706 -72660 73710 -71526
rect 73987 -71518 74064 -71517
rect 73987 -72652 73988 -71518
rect 74052 -72652 74064 -71518
rect 74360 -71537 74420 -71257
rect 74716 -71266 74720 -70084
rect 74796 -71266 74797 -70084
rect 75069 -71260 75070 -70078
rect 75146 -71260 75147 -70078
rect 75069 -71261 75147 -71260
rect 75427 -70078 75505 -70077
rect 75427 -71260 75428 -70078
rect 75504 -71260 75505 -70078
rect 75427 -71261 75505 -71260
rect 75781 -70078 75859 -70077
rect 75781 -71260 75782 -70078
rect 75858 -71260 75859 -70078
rect 75781 -71261 75859 -71260
rect 76135 -70078 76213 -70077
rect 76135 -71260 76136 -70078
rect 76212 -71260 76213 -70078
rect 76491 -71258 76492 -70076
rect 76568 -71258 76569 -70076
rect 76491 -71259 76569 -71258
rect 76852 -70087 76912 -70074
rect 77564 -70079 77624 -70078
rect 77197 -70080 77275 -70079
rect 76852 -70088 76931 -70087
rect 76135 -71261 76213 -71260
rect 74716 -71267 74797 -71266
rect 74716 -71529 74776 -71267
rect 73987 -72653 74064 -72652
rect 73641 -72661 73710 -72660
rect 73285 -72677 73354 -72676
rect 73294 -73704 73354 -72677
rect 73650 -73704 73710 -72661
rect 74004 -73704 74064 -72653
rect 74351 -71538 74420 -71537
rect 74351 -72672 74352 -71538
rect 74416 -72672 74420 -71538
rect 74713 -71530 74779 -71529
rect 74713 -72664 74714 -71530
rect 74778 -72664 74779 -71530
rect 75072 -71549 75132 -71261
rect 75428 -71537 75488 -71261
rect 75786 -71517 75846 -71261
rect 76140 -71517 76200 -71261
rect 76496 -71517 76556 -71259
rect 75763 -71518 75846 -71517
rect 75425 -71538 75491 -71537
rect 74713 -72665 74779 -72664
rect 75069 -71550 75135 -71549
rect 74351 -72673 74420 -72672
rect 74360 -73704 74420 -72673
rect 74716 -73704 74776 -72665
rect 75069 -72684 75070 -71550
rect 75134 -72684 75135 -71550
rect 75425 -72672 75426 -71538
rect 75490 -72672 75491 -71538
rect 75763 -72652 75764 -71518
rect 75828 -72652 75846 -71518
rect 75763 -72653 75846 -72652
rect 76127 -71518 76200 -71517
rect 76127 -72652 76128 -71518
rect 76192 -72652 76200 -71518
rect 76127 -72653 76200 -72652
rect 76477 -71518 76556 -71517
rect 76477 -72652 76478 -71518
rect 76542 -72652 76556 -71518
rect 76477 -72653 76556 -72652
rect 75425 -72673 75491 -72672
rect 75069 -72685 75135 -72684
rect 75072 -73704 75132 -72685
rect 75428 -73704 75488 -72673
rect 75786 -73704 75846 -72653
rect 76140 -73704 76200 -72653
rect 76496 -73704 76556 -72653
rect 76852 -71270 76854 -70088
rect 76930 -71270 76931 -70088
rect 77197 -71262 77198 -70080
rect 77274 -71262 77275 -70080
rect 77197 -71263 77275 -71262
rect 77553 -70080 77631 -70079
rect 77553 -71262 77554 -70080
rect 77630 -71262 77631 -70080
rect 77917 -71256 77918 -70074
rect 77994 -71256 77995 -70074
rect 79695 -70078 79773 -70077
rect 78276 -70083 78336 -70078
rect 78633 -70080 78711 -70079
rect 78991 -70080 79069 -70079
rect 77917 -71257 77995 -71256
rect 78271 -70084 78349 -70083
rect 77553 -71263 77631 -71262
rect 76852 -71271 76931 -71270
rect 76852 -71525 76912 -71271
rect 77210 -71525 77270 -71263
rect 76852 -71526 76919 -71525
rect 76852 -72660 76854 -71526
rect 76918 -72660 76919 -71526
rect 76852 -72661 76919 -72660
rect 77195 -71526 77270 -71525
rect 77195 -72660 77196 -71526
rect 77260 -72660 77270 -71526
rect 77564 -71537 77624 -71263
rect 77922 -71513 77982 -71257
rect 78271 -71266 78272 -70084
rect 78348 -71266 78349 -70084
rect 78633 -70086 78634 -70080
rect 78271 -71267 78349 -71266
rect 78632 -71262 78634 -70086
rect 78710 -71262 78711 -70080
rect 78632 -71263 78711 -71262
rect 78988 -71262 78992 -70080
rect 79068 -71262 79069 -70080
rect 78988 -71263 79069 -71262
rect 79344 -70083 79404 -70078
rect 79344 -70084 79423 -70083
rect 77195 -72661 77270 -72660
rect 76852 -73704 76912 -72661
rect 77210 -73704 77270 -72661
rect 77547 -71538 77624 -71537
rect 77547 -72672 77548 -71538
rect 77612 -72672 77624 -71538
rect 77909 -71514 77982 -71513
rect 77909 -72648 77910 -71514
rect 77974 -72648 77982 -71514
rect 78276 -71517 78336 -71267
rect 77909 -72649 77982 -72648
rect 77547 -72673 77624 -72672
rect 77564 -73704 77624 -72673
rect 77922 -73704 77982 -72649
rect 78273 -71518 78339 -71517
rect 78273 -72652 78274 -71518
rect 78338 -72652 78339 -71518
rect 78632 -71537 78692 -71263
rect 78273 -72653 78339 -72652
rect 78623 -71538 78692 -71537
rect 78276 -73704 78336 -72653
rect 78623 -72672 78624 -71538
rect 78688 -72672 78692 -71538
rect 78988 -71541 79048 -71263
rect 79344 -71266 79346 -70084
rect 79422 -71266 79423 -70084
rect 79695 -71260 79696 -70078
rect 79772 -71260 79773 -70078
rect 80058 -70083 80118 -70078
rect 80412 -70079 80472 -70078
rect 80768 -70079 80828 -70074
rect 81113 -70078 81191 -70077
rect 80411 -70080 80489 -70079
rect 79695 -71261 79773 -71260
rect 80051 -70084 80129 -70083
rect 79344 -71267 79423 -71266
rect 79344 -71517 79404 -71267
rect 79337 -71518 79404 -71517
rect 78623 -72673 78692 -72672
rect 78632 -73704 78692 -72673
rect 78987 -71542 79053 -71541
rect 78987 -72676 78988 -71542
rect 79052 -72676 79053 -71542
rect 79337 -72652 79338 -71518
rect 79402 -72652 79404 -71518
rect 79702 -71525 79762 -71261
rect 80051 -71266 80052 -70084
rect 80128 -71266 80129 -70084
rect 80411 -71262 80412 -70080
rect 80488 -71262 80489 -70080
rect 80411 -71263 80489 -71262
rect 80759 -70080 80837 -70079
rect 80759 -71262 80760 -70080
rect 80836 -71262 80837 -70080
rect 81113 -71260 81114 -70078
rect 81190 -71260 81191 -70078
rect 82194 -70079 82254 -70078
rect 81829 -70080 81907 -70079
rect 81482 -70083 81542 -70080
rect 81113 -71261 81191 -71260
rect 81477 -70084 81555 -70083
rect 80759 -71263 80837 -71262
rect 80051 -71267 80129 -71266
rect 79337 -72653 79404 -72652
rect 78987 -72677 79053 -72676
rect 78988 -73704 79048 -72677
rect 79344 -73704 79404 -72653
rect 79693 -71526 79762 -71525
rect 79693 -72660 79694 -71526
rect 79758 -72660 79762 -71526
rect 80058 -71529 80118 -71267
rect 79693 -72661 79762 -72660
rect 79702 -73704 79762 -72661
rect 80045 -71530 80118 -71529
rect 80045 -72664 80046 -71530
rect 80110 -72664 80118 -71530
rect 80412 -71537 80472 -71263
rect 80768 -71525 80828 -71263
rect 80045 -72665 80118 -72664
rect 80058 -73704 80118 -72665
rect 80399 -71538 80472 -71537
rect 80399 -72672 80400 -71538
rect 80464 -72672 80472 -71538
rect 80759 -71526 80828 -71525
rect 80759 -72660 80760 -71526
rect 80824 -72660 80828 -71526
rect 81124 -71537 81184 -71261
rect 81477 -71266 81478 -70084
rect 81554 -71266 81555 -70084
rect 81829 -71262 81830 -70080
rect 81906 -71262 81907 -70080
rect 81829 -71263 81907 -71262
rect 82175 -70080 82254 -70079
rect 82175 -71262 82176 -70080
rect 82252 -71262 82254 -70080
rect 82548 -70085 82608 -70080
rect 82906 -70083 82966 -70074
rect 83263 -70078 83264 -70070
rect 82893 -70084 82971 -70083
rect 82175 -71263 82254 -71262
rect 81477 -71267 81555 -71266
rect 81482 -71529 81542 -71267
rect 81838 -71529 81898 -71263
rect 81477 -71530 81543 -71529
rect 80759 -72661 80828 -72660
rect 80399 -72673 80472 -72672
rect 80412 -73704 80472 -72673
rect 80768 -73704 80828 -72661
rect 81121 -71538 81187 -71537
rect 81121 -72672 81122 -71538
rect 81186 -72672 81187 -71538
rect 81477 -72664 81478 -71530
rect 81542 -72664 81543 -71530
rect 81477 -72665 81543 -72664
rect 81838 -71530 81913 -71529
rect 81838 -72664 81848 -71530
rect 81912 -72664 81913 -71530
rect 82194 -71537 82254 -71263
rect 82533 -70086 82611 -70085
rect 82533 -71268 82534 -70086
rect 82610 -71268 82611 -70086
rect 82893 -71266 82894 -70084
rect 82970 -71266 82971 -70084
rect 82893 -71267 82971 -71266
rect 83262 -71252 83264 -70078
rect 83340 -71252 83341 -70070
rect 83262 -71253 83341 -71252
rect 83615 -70086 83693 -70085
rect 82533 -71269 82611 -71268
rect 81838 -72665 81913 -72664
rect 82183 -71538 82254 -71537
rect 81121 -72673 81187 -72672
rect 81124 -73704 81184 -72673
rect 81482 -73704 81542 -72665
rect 81838 -73704 81898 -72665
rect 82183 -72672 82184 -71538
rect 82248 -72672 82254 -71538
rect 82548 -71541 82608 -71269
rect 82183 -72673 82254 -72672
rect 82194 -73704 82254 -72673
rect 82541 -71542 82608 -71541
rect 82541 -72676 82542 -71542
rect 82606 -72676 82608 -71542
rect 82906 -71549 82966 -71267
rect 83262 -71529 83322 -71253
rect 83615 -71268 83616 -70086
rect 83692 -71268 83693 -70086
rect 83979 -70086 84057 -70085
rect 83979 -70088 83980 -70086
rect 83615 -71269 83693 -71268
rect 83974 -71268 83980 -70088
rect 84056 -71268 84057 -70086
rect 83974 -71269 84057 -71268
rect 83255 -71530 83322 -71529
rect 82541 -72677 82608 -72676
rect 82548 -73704 82608 -72677
rect 82905 -71550 82971 -71549
rect 82905 -72684 82906 -71550
rect 82970 -72684 82971 -71550
rect 83255 -72664 83256 -71530
rect 83320 -72664 83322 -71530
rect 83616 -71549 83676 -71269
rect 83974 -71529 84034 -71269
rect 83961 -71530 84034 -71529
rect 83255 -72665 83322 -72664
rect 82905 -72685 82971 -72684
rect 82906 -73704 82966 -72685
rect 83262 -73704 83322 -72665
rect 83611 -71550 83677 -71549
rect 83611 -72684 83612 -71550
rect 83676 -72684 83677 -71550
rect 83961 -72664 83962 -71530
rect 84026 -72664 84034 -71530
rect 83961 -72665 84034 -72664
rect 83611 -72685 83677 -72684
rect 83616 -73704 83676 -72685
rect 83974 -73704 84034 -72665
rect 68036 -74362 73354 -73704
rect 73568 -74354 78430 -73704
rect 67406 -84132 68036 -75561
rect 67406 -86766 68038 -84132
rect 69829 -84572 70489 -74362
rect 75616 -75636 76273 -74354
rect 78589 -74362 84068 -73704
rect 73390 -76775 74012 -75805
rect 73390 -79088 74006 -76775
rect 75616 -78968 76270 -75636
rect 73390 -80288 74022 -79088
rect 73390 -83626 74014 -80288
rect 75616 -80394 76273 -78968
rect 75616 -83860 76268 -80394
rect 79646 -83626 80270 -75864
rect 81770 -77206 82430 -74362
rect 81770 -77648 87454 -77206
rect 81770 -81902 82430 -77648
rect 87012 -81902 87454 -77648
rect 81770 -82335 87454 -81902
rect 81770 -82342 87438 -82335
rect 69832 -86516 70486 -84572
rect 75616 -86516 76273 -83860
rect 81770 -85477 82430 -82342
rect 84080 -82344 87438 -82342
rect 62934 -87632 64462 -87622
rect 60748 -87884 64462 -87632
rect 56240 -89338 59736 -89334
rect 56240 -89342 58674 -89338
rect 56240 -89346 56894 -89342
rect 56240 -90468 56534 -89346
rect 56610 -90464 56894 -89346
rect 56970 -89348 58674 -89342
rect 56970 -89350 58312 -89348
rect 56970 -89352 57956 -89350
rect 56970 -90464 57250 -89352
rect 56610 -90468 57250 -90464
rect 56240 -90474 57250 -90468
rect 57326 -90474 57600 -89352
rect 57676 -90472 57956 -89352
rect 58032 -90470 58312 -89350
rect 58388 -90460 58674 -89348
rect 58750 -89340 59736 -89338
rect 58750 -89350 59386 -89340
rect 58750 -90460 59024 -89350
rect 58388 -90470 59024 -90460
rect 58032 -90472 59024 -90470
rect 59100 -90462 59386 -89350
rect 59462 -90456 59736 -89340
rect 59812 -90456 60060 -89334
rect 59462 -90462 60060 -90456
rect 59100 -90472 60060 -90462
rect 57676 -90474 60060 -90472
rect 56240 -90682 60060 -90474
rect 60712 -89338 64462 -87884
rect 66760 -87398 68038 -86766
rect 68282 -87170 71916 -86516
rect 74146 -87170 77780 -86516
rect 81772 -86524 82429 -85477
rect 66760 -88642 67392 -87398
rect 68430 -87881 68490 -87170
rect 68430 -87882 68505 -87881
rect 60712 -89342 61676 -89338
rect 60712 -90464 60964 -89342
rect 61040 -89352 61676 -89342
rect 61040 -90464 61318 -89352
rect 60712 -90474 61318 -90464
rect 61394 -90460 61676 -89352
rect 61752 -89346 64462 -89338
rect 61752 -89348 63104 -89346
rect 61752 -90460 62036 -89348
rect 61394 -90470 62036 -90460
rect 62112 -89352 63104 -89348
rect 62112 -89354 62742 -89352
rect 62112 -90470 62392 -89354
rect 61394 -90474 62392 -90470
rect 60712 -90476 62392 -90474
rect 62468 -90474 62742 -89354
rect 62818 -90468 63104 -89352
rect 63180 -89360 63816 -89346
rect 63180 -90468 63458 -89360
rect 62818 -90474 63458 -90468
rect 62468 -90476 63458 -90474
rect 60712 -90482 63458 -90476
rect 63534 -90468 63816 -89360
rect 63892 -89352 64462 -89346
rect 63892 -90468 64176 -89352
rect 63534 -90474 64176 -90468
rect 64252 -90474 64462 -89352
rect 68430 -89014 68436 -87882
rect 68504 -89014 68505 -87882
rect 68430 -89015 68505 -89014
rect 68786 -87889 68846 -87170
rect 69142 -87889 69202 -87170
rect 68786 -87890 68867 -87889
rect 68430 -89307 68490 -89015
rect 68786 -89022 68798 -87890
rect 68866 -89022 68867 -87890
rect 68786 -89023 68867 -89022
rect 69142 -87890 69217 -87889
rect 69142 -89022 69148 -87890
rect 69216 -89022 69217 -87890
rect 69142 -89023 69217 -89022
rect 69498 -87891 69558 -87170
rect 69854 -87887 69914 -87170
rect 69854 -87888 69929 -87887
rect 69498 -87892 69575 -87891
rect 68786 -89307 68846 -89023
rect 69142 -89307 69202 -89023
rect 69498 -89024 69506 -87892
rect 69574 -89024 69575 -87892
rect 69498 -89025 69575 -89024
rect 69854 -89020 69860 -87888
rect 69928 -89020 69929 -87888
rect 69854 -89021 69929 -89020
rect 70210 -87893 70270 -87170
rect 70566 -87889 70626 -87170
rect 70566 -87890 70643 -87889
rect 70210 -87894 70281 -87893
rect 68430 -89308 68509 -89307
rect 68430 -90440 68440 -89308
rect 68508 -90440 68509 -89308
rect 68430 -90441 68509 -90440
rect 68786 -89308 68865 -89307
rect 68786 -90440 68796 -89308
rect 68864 -90440 68865 -89308
rect 68786 -90441 68865 -90440
rect 69142 -89308 69219 -89307
rect 69142 -90440 69150 -89308
rect 69218 -90440 69219 -89308
rect 69142 -90441 69219 -90440
rect 69498 -89309 69558 -89025
rect 69498 -89310 69569 -89309
rect 68430 -90466 68490 -90441
rect 68786 -90468 68846 -90441
rect 69142 -90456 69202 -90441
rect 69498 -90442 69500 -89310
rect 69568 -90442 69569 -89310
rect 69499 -90443 69569 -90442
rect 69854 -89315 69914 -89021
rect 70210 -89026 70212 -87894
rect 70280 -89026 70281 -87894
rect 70210 -89027 70281 -89026
rect 70566 -89022 70574 -87890
rect 70642 -89022 70643 -87890
rect 70566 -89023 70643 -89022
rect 70924 -87893 70984 -87170
rect 70924 -87894 70997 -87893
rect 70210 -89315 70270 -89027
rect 70566 -89313 70626 -89023
rect 70924 -89026 70928 -87894
rect 70996 -89026 70997 -87894
rect 70924 -89027 70997 -89026
rect 71278 -87897 71338 -87170
rect 71636 -87893 71696 -87170
rect 74320 -87879 74380 -87170
rect 74320 -87880 74401 -87879
rect 71636 -87894 71713 -87893
rect 71278 -87898 71355 -87897
rect 70924 -89311 70984 -89027
rect 71278 -89030 71286 -87898
rect 71354 -89030 71355 -87898
rect 71278 -89031 71355 -89030
rect 71636 -89026 71644 -87894
rect 71712 -89026 71713 -87894
rect 71636 -89027 71713 -89026
rect 74320 -89012 74332 -87880
rect 74400 -89012 74401 -87880
rect 74320 -89013 74401 -89012
rect 74676 -87887 74736 -87170
rect 75032 -87887 75092 -87170
rect 74676 -87888 74763 -87887
rect 70924 -89312 70995 -89311
rect 70566 -89314 70639 -89313
rect 69854 -89316 69925 -89315
rect 69854 -90448 69856 -89316
rect 69924 -90448 69925 -89316
rect 70210 -89316 70289 -89315
rect 70210 -90432 70220 -89316
rect 69854 -90449 69925 -90448
rect 70219 -90448 70220 -90432
rect 70288 -90448 70289 -89316
rect 70219 -90449 70289 -90448
rect 70566 -90446 70570 -89314
rect 70638 -90446 70639 -89314
rect 70924 -90442 70926 -89312
rect 70925 -90444 70926 -90442
rect 70994 -90444 70995 -89312
rect 70925 -90445 70995 -90444
rect 71278 -89315 71338 -89031
rect 71636 -89315 71696 -89027
rect 74320 -89305 74380 -89013
rect 74676 -89020 74694 -87888
rect 74762 -89020 74763 -87888
rect 74676 -89021 74763 -89020
rect 75032 -87888 75113 -87887
rect 75032 -89020 75044 -87888
rect 75112 -89020 75113 -87888
rect 75032 -89021 75113 -89020
rect 75388 -87889 75448 -87170
rect 75744 -87885 75804 -87170
rect 75744 -87886 75825 -87885
rect 75388 -87890 75471 -87889
rect 74676 -89305 74736 -89021
rect 75032 -89305 75092 -89021
rect 75388 -89022 75402 -87890
rect 75470 -89022 75471 -87890
rect 75388 -89023 75471 -89022
rect 75744 -89018 75756 -87886
rect 75824 -89018 75825 -87886
rect 75744 -89019 75825 -89018
rect 76100 -87891 76160 -87170
rect 76456 -87887 76516 -87170
rect 76456 -87888 76539 -87887
rect 76100 -87892 76177 -87891
rect 74320 -89306 74405 -89305
rect 71278 -89316 71355 -89315
rect 70566 -90447 70639 -90446
rect 69854 -90456 69914 -90449
rect 70566 -90458 70626 -90447
rect 71278 -90448 71286 -89316
rect 71354 -90448 71355 -89316
rect 71278 -90449 71355 -90448
rect 71633 -89316 71703 -89315
rect 71633 -90448 71634 -89316
rect 71702 -90448 71703 -89316
rect 71633 -90449 71703 -90448
rect 74320 -90438 74336 -89306
rect 74404 -90438 74405 -89306
rect 74320 -90439 74405 -90438
rect 74676 -89306 74761 -89305
rect 74676 -90438 74692 -89306
rect 74760 -90438 74761 -89306
rect 74676 -90439 74761 -90438
rect 75032 -89306 75115 -89305
rect 75032 -90438 75046 -89306
rect 75114 -90438 75115 -89306
rect 75032 -90439 75115 -90438
rect 75388 -89307 75448 -89023
rect 75388 -89308 75465 -89307
rect 71278 -90456 71338 -90449
rect 74320 -90468 74380 -90439
rect 74676 -90460 74736 -90439
rect 75032 -90450 75092 -90439
rect 75388 -90440 75396 -89308
rect 75464 -90440 75465 -89308
rect 75388 -90441 75465 -90440
rect 75744 -89313 75804 -89019
rect 76100 -89024 76108 -87892
rect 76176 -89024 76177 -87892
rect 76100 -89025 76177 -89024
rect 76456 -89020 76470 -87888
rect 76538 -89020 76539 -87888
rect 76456 -89021 76539 -89020
rect 76814 -87891 76874 -87170
rect 76814 -87892 76893 -87891
rect 76100 -89313 76160 -89025
rect 76456 -89311 76516 -89021
rect 76814 -89024 76824 -87892
rect 76892 -89024 76893 -87892
rect 76814 -89025 76893 -89024
rect 77168 -87895 77228 -87170
rect 77526 -87891 77586 -87170
rect 80288 -87172 83922 -86524
rect 80450 -87873 80510 -87172
rect 80445 -87874 80515 -87873
rect 77526 -87892 77609 -87891
rect 77168 -87896 77251 -87895
rect 76814 -89309 76874 -89025
rect 77168 -89028 77182 -87896
rect 77250 -89028 77251 -87896
rect 77168 -89029 77251 -89028
rect 77526 -89024 77540 -87892
rect 77608 -89024 77609 -87892
rect 80445 -89006 80446 -87874
rect 80514 -89006 80515 -87874
rect 80445 -89007 80515 -89006
rect 80806 -87881 80866 -87172
rect 81162 -87881 81222 -87172
rect 80806 -87882 80877 -87881
rect 77526 -89025 77609 -89024
rect 76814 -89310 76891 -89309
rect 76456 -89312 76535 -89311
rect 75744 -89314 75821 -89313
rect 75388 -90460 75448 -90441
rect 75744 -90446 75752 -89314
rect 75820 -90446 75821 -89314
rect 75751 -90447 75821 -90446
rect 76100 -89314 76185 -89313
rect 76100 -90446 76116 -89314
rect 76184 -90446 76185 -89314
rect 76456 -90444 76466 -89312
rect 76534 -90444 76535 -89312
rect 76456 -90445 76535 -90444
rect 76814 -90442 76822 -89310
rect 76890 -90442 76891 -89310
rect 77168 -89313 77228 -89029
rect 77526 -89313 77586 -89025
rect 80450 -89299 80510 -89007
rect 80806 -89014 80808 -87882
rect 80876 -89014 80877 -87882
rect 80806 -89015 80877 -89014
rect 81157 -87882 81227 -87881
rect 81157 -89014 81158 -87882
rect 81226 -89014 81227 -87882
rect 81518 -87883 81578 -87172
rect 81874 -87879 81934 -87172
rect 81869 -87880 81939 -87879
rect 81157 -89015 81227 -89014
rect 81515 -87884 81585 -87883
rect 80806 -89299 80866 -89015
rect 81162 -89299 81222 -89015
rect 81515 -89016 81516 -87884
rect 81584 -89016 81585 -87884
rect 81869 -89012 81870 -87880
rect 81938 -89012 81939 -87880
rect 82230 -87885 82290 -87172
rect 82586 -87881 82646 -87172
rect 82583 -87882 82653 -87881
rect 81869 -89013 81939 -89012
rect 82221 -87886 82291 -87885
rect 81515 -89017 81585 -89016
rect 80449 -89300 80519 -89299
rect 77168 -89314 77251 -89313
rect 77168 -90436 77182 -89314
rect 76814 -90443 76891 -90442
rect 76456 -90446 76516 -90445
rect 76100 -90447 76185 -90446
rect 76100 -90450 76160 -90447
rect 76814 -90460 76874 -90443
rect 77181 -90446 77182 -90436
rect 77250 -90446 77251 -89314
rect 77526 -89314 77599 -89313
rect 77526 -90446 77530 -89314
rect 77598 -90446 77599 -89314
rect 80449 -90432 80450 -89300
rect 80518 -90432 80519 -89300
rect 80449 -90433 80519 -90432
rect 80805 -89300 80875 -89299
rect 80805 -90432 80806 -89300
rect 80874 -90432 80875 -89300
rect 80805 -90433 80875 -90432
rect 81159 -89300 81229 -89299
rect 81159 -90432 81160 -89300
rect 81228 -90432 81229 -89300
rect 81518 -89301 81578 -89017
rect 81159 -90433 81229 -90432
rect 81509 -89302 81579 -89301
rect 80450 -90436 80510 -90433
rect 80806 -90446 80866 -90433
rect 81162 -90436 81222 -90433
rect 81509 -90434 81510 -89302
rect 81578 -90434 81579 -89302
rect 81874 -89307 81934 -89013
rect 82221 -89018 82222 -87886
rect 82290 -89018 82291 -87886
rect 82583 -89014 82584 -87882
rect 82652 -89014 82653 -87882
rect 82944 -87885 83004 -87172
rect 82583 -89015 82653 -89014
rect 82937 -87886 83007 -87885
rect 82221 -89019 82291 -89018
rect 82230 -89307 82290 -89019
rect 82586 -89305 82646 -89015
rect 82937 -89018 82938 -87886
rect 83006 -89018 83007 -87886
rect 83298 -87889 83358 -87172
rect 83656 -87885 83716 -87172
rect 83653 -87886 83723 -87885
rect 82937 -89019 83007 -89018
rect 83295 -87890 83365 -87889
rect 82944 -89303 83004 -89019
rect 83295 -89022 83296 -87890
rect 83364 -89022 83365 -87890
rect 83653 -89018 83654 -87886
rect 83722 -89018 83723 -87886
rect 83653 -89019 83723 -89018
rect 83295 -89023 83365 -89022
rect 82935 -89304 83005 -89303
rect 82579 -89306 82649 -89305
rect 81509 -90435 81579 -90434
rect 81865 -89308 81935 -89307
rect 81518 -90446 81578 -90435
rect 81865 -90440 81866 -89308
rect 81934 -90440 81935 -89308
rect 81865 -90441 81935 -90440
rect 82229 -89308 82299 -89307
rect 82229 -90440 82230 -89308
rect 82298 -90440 82299 -89308
rect 82579 -90438 82580 -89306
rect 82648 -90438 82649 -89306
rect 82935 -90436 82936 -89304
rect 83004 -90436 83005 -89304
rect 83298 -89307 83358 -89023
rect 83656 -89307 83716 -89019
rect 82935 -90437 83005 -90436
rect 83295 -89308 83365 -89307
rect 82579 -90439 82649 -90438
rect 82229 -90441 82299 -90440
rect 77181 -90447 77251 -90446
rect 77529 -90447 77599 -90446
rect 81874 -90450 81934 -90441
rect 82230 -90446 82290 -90441
rect 82586 -90450 82646 -90439
rect 82944 -90450 83004 -90437
rect 83295 -90440 83296 -89308
rect 83364 -90440 83365 -89308
rect 83295 -90441 83365 -90440
rect 83643 -89308 83716 -89307
rect 83643 -90440 83644 -89308
rect 83712 -90440 83716 -89308
rect 83643 -90441 83716 -90440
rect 83298 -90450 83358 -90441
rect 83656 -90446 83716 -90441
rect 63534 -90482 64462 -90474
rect 60712 -90680 64462 -90482
rect 60712 -90682 63412 -90680
rect 60712 -90686 62172 -90682
use sky130_fd_pr__nfet_01v8_X8JY7K  sky130_fd_pr__nfet_01v8_X8JY7K_0
timestamp 1607735006
transform 1 0 58169 0 1 -89898
box -1947 -810 1947 810
use sky130_fd_pr__nfet_01v8_X8JY7K  sky130_fd_pr__nfet_01v8_X8JY7K_1
timestamp 1607735006
transform 1 0 62605 0 1 -89896
box -1947 -810 1947 810
use via_m2_m3  via_m2_m3_1
array 0 9 84 0 9 84
timestamp 1606703199
transform 1 0 54904 0 1 -89644
box -14 -14 70 70
use via_m2_m3  via_m2_m3_2
array 0 9 84 0 9 84
timestamp 1606703199
transform 1 0 54908 0 1 -90588
box -14 -14 70 70
use via_li_m1  via_li_m1_0
array 0 7 72 0 19 74
timestamp 1606675505
transform 1 0 64650 0 1 -90538
box 4 0 76 74
use via_m3_m4  via_m3_m4_12
array 0 9 104 0 5 104
timestamp 1606691473
transform 1 0 64242 0 1 -92090
box -20 -20 84 84
use sky130_fd_pr__nfet_01v8_XGTW7K  sky130_fd_pr__nfet_01v8_XGTW7K_0
timestamp 1607714484
transform 1 0 70073 0 1 -89151
box -1947 -1519 1947 1519
use via_m2_m3  via_m2_m3_9
array 0 24 84 0 7 84
timestamp 1606703199
transform 1 0 65434 0 1 -90500
box -14 -14 70 70
use via_li_m1  via_li_m1_4
array 0 125 72 0 4 74
timestamp 1606675505
transform 1 0 56266 0 1 -89016
box 4 0 76 74
use via_li_m1  via_li_m1_11
array 0 19 72 0 34 74
timestamp 1606675505
transform 1 0 78208 0 1 -90402
box 4 0 76 74
use via_li_m1  via_li_m1_10
array 0 19 72 0 34 74
timestamp 1606675505
transform 1 0 72256 0 1 -90430
box 4 0 76 74
use sky130_fd_pr__nfet_01v8_XGTW7K  sky130_fd_pr__nfet_01v8_XGTW7K_2
timestamp 1607714484
transform 1 0 82085 0 1 -89151
box -1947 -1519 1947 1519
use sky130_fd_pr__nfet_01v8_XGTW7K  sky130_fd_pr__nfet_01v8_XGTW7K_1
timestamp 1607714484
transform 1 0 75961 0 1 -89151
box -1947 -1519 1947 1519
use via_li_m1  via_li_m1_12
array 0 19 72 0 34 74
timestamp 1606675505
transform 1 0 84378 0 1 -90444
box 4 0 76 74
use via_m2_m3  via_m2_m3_0
array 0 369 84 0 9 84
timestamp 1606703199
transform 1 0 55070 0 1 -91866
box -14 -14 70 70
use via_li_m1  via_li_m1_5
array 0 429 72 0 9 74
timestamp 1606675505
transform 1 0 55060 0 1 -91886
box 4 0 76 74
use via_m3_m4  via_m3_m4_1
array 0 5 104 0 3 104
timestamp 1606691473
transform 1 0 65926 0 1 -87360
box -20 -20 84 84
use via_m3_m4  via_m3_m4_6
array 0 29 104 0 5 104
timestamp 1606691473
transform 1 0 74236 0 1 -87124
box -20 -20 84 84
use via_m3_m4  via_m3_m4_7
array 0 29 104 0 5 104
timestamp 1606691473
transform 1 0 68356 0 1 -87124
box -20 -20 84 84
use via_m3_m4  via_m3_m4_5
array 0 29 104 0 5 104
timestamp 1606691473
transform 1 0 80434 0 1 -87124
box -20 -20 84 84
use via_m2_m3  via_m2_m3_7
array 0 5 84 0 3 84
timestamp 1606703199
transform 1 0 65948 0 1 -87378
box -14 -14 70 70
use sky130_fd_pr__pfet_01v8_JXF9S2  sky130_fd_pr__pfet_01v8_JXF9S2_3
timestamp 1607731921
transform 1 0 60320 0 1 -86353
box -4172 -1537 4172 1537
use via_m3_m4  via_m3_m4_11
array 0 5 104 0 3 104
timestamp 1606691473
transform 1 0 66732 0 1 -88584
box -20 -20 84 84
use sky130_fd_pr__cap_mim_m3_1_BLS9H9  sky130_fd_pr__cap_mim_m3_1_BLS9H9_4
timestamp 1606520558
transform -1 0 69939 0 1 -82050
box -1941 -1600 1941 1600
use sky130_fd_pr__cap_mim_m3_1_BLS9H9  sky130_fd_pr__cap_mim_m3_1_BLS9H9_1
timestamp 1606520558
transform -1 0 75899 0 1 -82032
box -1941 -1600 1941 1600
use sky130_fd_pr__cap_mim_m3_1_BLS9H9  sky130_fd_pr__cap_mim_m3_1_BLS9H9_3
timestamp 1606520558
transform -1 0 82189 0 1 -82052
box -1941 -1600 1941 1600
use sky130_fd_pr__pfet_01v8_JXF9S2  sky130_fd_pr__pfet_01v8_JXF9S2_2
timestamp 1607731921
transform 1 0 60344 0 1 -82535
box -4172 -1537 4172 1537
use via_li_m1  via_li_m1_6
array 0 109 72 0 2 74
timestamp 1606675505
transform 1 0 56292 0 1 -84564
box 4 0 76 74
use via_m3_m4  via_m3_m4_8
array 0 3 104 0 5 104
timestamp 1606691473
transform 1 0 79708 0 1 -79968
box -20 -20 84 84
use sky130_fd_pr__cap_mim_m3_1_BLS9H9  sky130_fd_pr__cap_mim_m3_1_BLS9H9_0
timestamp 1606520558
transform -1 0 75933 0 1 -77394
box -1941 -1600 1941 1600
use sky130_fd_pr__cap_mim_m3_1_BLS9H9  sky130_fd_pr__cap_mim_m3_1_BLS9H9_2
timestamp 1606520558
transform -1 0 82189 0 1 -77554
box -1941 -1600 1941 1600
use sky130_fd_pr__cap_mim_m3_1_BLS9H9  sky130_fd_pr__cap_mim_m3_1_BLS9H9_5
timestamp 1606520558
transform -1 0 69957 0 1 -77200
box -1941 -1600 1941 1600
use via_m3_m4  via_m3_m4_10
array 0 3 104 0 5 104
timestamp 1606691473
transform 1 0 67502 0 1 -79996
box -20 -20 84 84
use via_m3_m4  via_m3_m4_9
array 0 3 104 0 5 104
timestamp 1606691473
transform 1 0 73448 0 1 -79996
box -20 -20 84 84
use sky130_fd_pr__pfet_01v8_JXF9S2  sky130_fd_pr__pfet_01v8_JXF9S2_1
timestamp 1607731921
transform 1 0 60342 0 1 -78567
box -4172 -1537 4172 1537
use via_li_m1  via_li_m1_7
array 0 109 72 0 2 74
timestamp 1606675505
transform 1 0 56298 0 1 -80712
box 4 0 76 74
use via_li_m1  via_li_m1_8
array 0 109 72 0 2 74
timestamp 1606675505
transform 1 0 56292 0 1 -76728
box 4 0 76 74
use via_m3_m4  via_m3_m4_4
array 0 44 104 0 5 104
timestamp 1606691473
transform 1 0 78666 0 1 -74318
box -20 -20 84 84
use via_m3_m4  via_m3_m4_2
array 0 44 104 0 5 104
timestamp 1606691473
transform 1 0 68276 0 1 -74326
box -20 -20 84 84
use via_m3_m4  via_m3_m4_3
array 0 44 104 0 5 104
timestamp 1606691473
transform 1 0 73654 0 1 -74332
box -20 -20 84 84
use sky130_fd_pr__pfet_01v8_JXF9S2  sky130_fd_pr__pfet_01v8_JXF9S2_0
timestamp 1607731921
transform 1 0 60350 0 1 -74719
box -4172 -1537 4172 1537
use via_li_m1  via_li_m1_13
array 0 19 72 0 34 74
timestamp 1606675505
transform 1 0 84582 0 1 -72614
box 4 0 76 74
use via_m2_m3  via_m2_m3_8
array 0 99 84 0 5 84
timestamp 1606703199
transform 1 0 56326 0 1 -73104
box -14 -14 70 70
use sky130_fd_pr__pfet_01v8_VXT95W  sky130_fd_pr__pfet_01v8_VXT95W_1
timestamp 1607649912
transform 1 0 76169 0 1 -71413
box -8177 -1537 8177 1537
use sky130_fd_pr__pfet_01v8_VXTF3X  sky130_fd_pr__pfet_01v8_VXTF3X_1
timestamp 1608072956
transform 1 0 62583 0 1 -70705
box -1947 -819 1947 819
use sky130_fd_pr__pfet_01v8_VXTQ3X  sky130_fd_pr__pfet_01v8_VXTQ3X_1
timestamp 1608072348
transform 1 0 57913 0 1 -70707
box -1769 -819 1769 819
use via_li_m1  via_li_m1_9
array 0 109 72 0 2 74
timestamp 1606675505
transform 1 0 56320 0 1 -73122
box 4 0 76 74
use via_m2_m3  via_m2_m3_3
array 0 99 84 0 3 84
timestamp 1606703199
transform 1 0 56158 0 1 -69674
box -14 -14 70 70
use via_li_m1  via_li_m1_1
array 0 119 72 0 3 74
timestamp 1606675505
transform 1 0 56146 0 1 -69710
box 4 0 76 74
use via_m2_m3  via_m2_m3_6
array 0 5 84 0 3 84
timestamp 1606703199
transform 1 0 65940 0 1 -69690
box -14 -14 70 70
use via_m3_m4  via_m3_m4_0
array 0 5 104 0 3 104
timestamp 1606691473
transform 1 0 65968 0 1 -69752
box -20 -20 84 84
use via_m2_m3  via_m2_m3_4
array 0 99 84 0 3 84
timestamp 1606703199
transform 1 0 68044 0 1 -69644
box -14 -14 70 70
use via_li_m1  via_li_m1_3
array 0 199 72 0 3 74
timestamp 1606675505
transform 1 0 69014 0 1 -69672
box 4 0 76 74
use via_m2_m3  via_m2_m3_5
array 0 99 84 0 3 84
timestamp 1606703199
transform 1 0 76440 0 1 -69640
box -14 -14 70 70
use sky130_fd_pr__nfet_01v8_PGN2UQ  sky130_fd_pr__nfet_01v8_PGN2UQ_0
timestamp 1608096578
transform 1 0 66705 0 1 -88335
box -10253 -937 701 18252
use via_li_m1  via_li_m1_2
array 0 219 -72 0 3 74
timestamp 1606675505
transform 0 1 55742 -1 0 -88278
box 4 0 76 74
<< labels >>
rlabel metal4 87012 -82335 87454 -77206 1 vout
rlabel metal2 53804 -76772 54966 -76432 1 vin_n
rlabel metal2 53796 -84634 54958 -84294 1 vin_p
rlabel metal3 56230 -73064 65354 -72630 1 vp
rlabel metal2 52320 -69842 52878 -69270 1 vdd
rlabel metal2 52394 -71478 52800 -71338 1 iref
rlabel metal2 59910 -89258 60874 -89126 1 vbn
rlabel metal2 54869 -91946 56021 -91031 1 vss
<< end >>
