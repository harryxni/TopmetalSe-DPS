magic
tech sky130B
magscale 1 2
timestamp 1662069552
<< metal1 >>
rect -80 3120 4925 3270
rect 5075 3120 5081 3270
rect 3490 1590 5850 1650
rect 5910 1590 5916 1650
rect 90 330 420 480
rect 3085 330 3585 480
rect 3735 330 4280 480
<< via1 >>
rect 4925 3120 5075 3270
rect 5850 1590 5910 1650
rect 3585 330 3735 480
<< metal2 >>
rect 4379 738 4542 3611
rect 4925 3270 5075 3276
rect 4916 3120 4925 3270
rect 5075 3120 5084 3270
rect 4925 3114 5075 3120
rect 4379 682 4432 738
rect 4488 682 4542 738
rect 3585 480 3735 486
rect 3576 330 3585 480
rect 3735 330 3744 480
rect 3585 324 3735 330
rect 4379 -231 4542 682
rect 5375 2098 5585 3645
rect 5375 2042 5452 2098
rect 5508 2042 5585 2098
rect 5375 -255 5585 2042
rect 5850 1650 5910 1659
rect 5850 1581 5910 1590
<< via2 >>
rect 4925 3120 5075 3270
rect 4432 682 4488 738
rect 3585 330 3735 480
rect 5452 2042 5508 2098
rect 5850 1590 5910 1650
<< metal3 >>
rect 4920 3270 4930 3275
rect 4920 3120 4925 3270
rect 4920 3115 4930 3120
rect 5080 3115 5086 3275
rect -80 2990 250 3050
rect -80 2790 60 2850
rect -80 2490 160 2550
rect 6608 2232 6672 2238
rect 3500 2170 6608 2230
rect 6608 2162 6672 2168
rect 5447 2100 5513 2103
rect 3470 2098 5513 2100
rect 3470 2042 5452 2098
rect 5508 2042 5513 2098
rect 3470 2040 5513 2042
rect 5447 2037 5513 2040
rect 6168 1932 6232 1938
rect 3500 1870 6168 1930
rect 6168 1862 6232 1868
rect 5820 1655 5930 1680
rect 5820 1591 5845 1655
rect 5915 1591 5930 1655
rect 5820 1590 5850 1591
rect 5910 1590 5930 1591
rect 5820 1560 5930 1590
rect 4427 740 4493 743
rect -80 680 80 740
rect 3470 738 4493 740
rect 3470 682 4432 738
rect 4488 682 4493 738
rect 3470 680 4493 682
rect 4427 677 4493 680
rect 3470 485 3780 490
rect 3470 480 3590 485
rect 3470 330 3585 480
rect 3470 325 3590 330
rect 3740 325 3780 485
rect 3470 310 3780 325
rect 3940 480 4090 486
rect 4090 330 4280 480
rect 3940 324 4090 330
<< via3 >>
rect 4930 3270 5080 3275
rect 4930 3120 5075 3270
rect 5075 3120 5080 3270
rect 4930 3115 5080 3120
rect 6608 2168 6672 2232
rect 6168 1868 6232 1932
rect 5845 1650 5915 1655
rect 5845 1591 5850 1650
rect 5850 1591 5910 1650
rect 5910 1591 5915 1650
rect 3590 480 3740 485
rect 3590 330 3735 480
rect 3735 330 3740 480
rect 3590 325 3740 330
rect 3940 330 4090 480
<< metal4 >>
rect 3805 3160 4195 3640
rect 4800 3490 5200 3650
rect 4800 3355 4855 3490
rect 5175 3370 5200 3490
rect 5175 3355 5210 3370
rect 3835 3030 4185 3160
rect 4800 3035 4850 3355
rect 5180 3035 5210 3355
rect 3589 485 3741 486
rect 3589 325 3590 485
rect 3740 480 3741 485
rect 4800 2820 4855 3035
rect 5175 3030 5210 3035
rect 5175 2820 5200 3030
rect 5850 1656 5910 3640
rect 6170 1933 6230 3640
rect 6460 3455 6840 3560
rect 6460 2360 6500 3455
rect 6460 2040 6480 2360
rect 6167 1932 6233 1933
rect 6167 1868 6168 1932
rect 6232 1868 6233 1932
rect 6167 1867 6233 1868
rect 5844 1655 5916 1656
rect 5844 1591 5845 1655
rect 5915 1591 5916 1655
rect 5844 1590 5916 1591
rect 3740 330 3855 480
rect 4175 330 4230 480
rect 3740 325 3741 330
rect 3589 324 3741 325
rect 4830 110 5190 290
rect 5850 -220 5910 1590
rect 6170 -270 6230 1867
rect 6460 570 6500 2040
rect 6810 570 6840 3455
rect 6460 -310 6840 570
<< via4 >>
rect 4855 3355 5175 3490
rect 4850 3275 5180 3355
rect 4850 3115 4930 3275
rect 4930 3115 5080 3275
rect 5080 3115 5180 3275
rect 4850 3035 5180 3115
rect 3855 480 4175 3030
rect 4855 650 5175 3035
rect 6500 2360 6810 3455
rect 6480 2232 6810 2360
rect 6480 2168 6608 2232
rect 6608 2168 6672 2232
rect 6672 2168 6810 2232
rect 6480 2040 6810 2168
rect 3855 330 3940 480
rect 3940 330 4090 480
rect 4090 330 4175 480
rect 3855 170 4175 330
rect 6500 570 6810 2040
<< metal5 >>
rect 3805 3320 4195 3640
rect 4800 3490 5200 3650
rect 4800 3355 4855 3490
rect 5175 3379 5200 3490
rect 6460 3455 6840 3630
rect 5175 3355 5213 3379
rect 3805 3030 4205 3320
rect 3805 170 3855 3030
rect 4175 170 4205 3030
rect 4800 3035 4850 3355
rect 5180 3035 5213 3355
rect 4800 2820 4855 3035
rect 3805 -120 4205 170
rect 4805 650 4855 2820
rect 5175 3011 5213 3035
rect 5175 650 5205 3011
rect 6460 2384 6500 3455
rect 6456 2360 6500 2384
rect 6456 2040 6480 2360
rect 6456 2016 6500 2040
rect 4805 -120 5205 650
rect 6460 570 6500 2016
rect 6810 570 6840 3455
rect 6460 -310 6840 570
use pixel  pixel_0
timestamp 1662068818
transform 1 0 470 0 1 3000
box -470 -3000 3090 570
<< end >>
