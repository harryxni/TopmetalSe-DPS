magic
tech sky130B
timestamp 1662181890
use bottom_left_pixel  bottom_left_pixel_0
timestamp 1662181890
transform 1 0 1410 0 1 -3000
box -1410 -2245 1975 1820
use bottom_pixel  bottom_pixel_0
timestamp 1662180122
transform 1 0 3145 0 1 -1535
box -385 -3710 1740 320
use bottom_right_pixel  bottom_right_pixel_0
timestamp 1662181774
transform 1 0 4645 0 1 -1535
box -385 -3710 3185 360
use left_pixel  left_pixel_0
timestamp 1662181890
transform 1 0 1410 0 1 -1500
box -1410 -65 1780 1820
use pixel  pixel_0
timestamp 1662180122
transform 1 0 3145 0 1 0
box -235 -1500 1545 285
use right_pixel  right_pixel_0
timestamp 1662181774
transform 1 0 4410 0 1 -1500
box -40 -155 3420 1825
use top_left_pixel  top_left_pixel_0
timestamp 1662180174
transform 1 0 1410 0 1 75
box -1410 -75 1785 2190
use top_pixel  top_pixel_0
timestamp 1662180122
transform 1 0 2915 0 1 75
box -5 0 1780 2190
use top_right_pixel  top_right_pixel_0
timestamp 1662181890
transform 1 0 4410 0 1 75
box -40 -155 3420 2190
<< end >>
