magic
tech sky130B
magscale 1 2
timestamp 1662181890
<< locali >>
rect 53780 204191 53850 204462
<< viali >>
rect 53780 204462 53850 204532
<< metal1 >>
rect 24140 692850 26600 692870
rect 22490 692780 26600 692850
rect 22490 691070 22560 692780
rect 26520 691070 26600 692780
rect 22490 690940 26600 691070
rect 24140 690410 26600 690940
rect 26190 689470 39770 689570
rect 26190 688990 36060 689470
rect 26200 687790 36060 688990
rect 39510 689460 39770 689470
rect 39510 687790 42700 689460
rect 26200 687620 42700 687790
rect 26663 683632 27687 687620
rect 29716 683675 30585 687620
rect 31111 683649 31609 687620
rect 36390 686900 42700 687620
rect 31111 683145 31609 683151
rect 29716 682800 30585 682806
rect 26663 682322 27687 682328
rect 57310 224245 57316 226314
rect 59385 224245 59391 226314
rect 57316 221685 59385 224245
rect 18576 219616 59385 221685
rect 18576 160435 20645 219616
rect 57316 219526 59385 219616
rect 53715 205825 59960 206575
rect 44080 204950 46260 205280
rect 53879 204990 53991 205825
rect 54079 204990 54191 205825
rect 54279 204990 54391 205825
rect 54479 204990 54591 205825
rect 54679 204990 54791 205825
rect 54879 204990 54991 205825
rect 55079 204990 55191 205825
rect 55279 204990 55391 205825
rect 55479 204990 55591 205825
rect 55679 204990 55791 205825
rect 59210 204990 59960 205825
rect 545850 205030 549270 205460
rect 60625 204990 549270 205030
rect 44080 201770 44290 204950
rect 46040 203890 46260 204950
rect 53720 204960 549270 204990
rect 53720 204930 60690 204960
rect 53720 204740 55880 204930
rect 57195 204740 60690 204930
rect 53720 204700 60690 204740
rect 53768 204456 53774 204538
rect 53844 204532 53862 204538
rect 53850 204462 53862 204532
rect 53844 204456 53862 204462
rect 49580 204410 49640 204416
rect 49640 204350 53720 204410
rect 49580 204344 49640 204350
rect 53660 204120 53720 204350
rect 53520 203905 53610 204120
rect 53405 203890 53765 203905
rect 46040 203870 53765 203890
rect 53490 203835 53765 203870
rect 53490 203645 53680 203835
rect 53490 203470 53685 203645
rect 46040 203370 53685 203470
rect 46040 203360 53630 203370
rect 46040 203342 53670 203360
rect 46040 203297 53685 203342
rect 46040 203170 53580 203297
rect 56375 203170 57125 204700
rect 58105 203170 58855 204700
rect 59210 203170 59960 204700
rect 60625 203170 60690 204700
rect 46040 202800 46260 203170
rect 52270 202800 52570 203170
rect 46040 202500 52570 202800
rect 56225 202620 60690 203170
rect 46040 202040 46260 202500
rect 52270 202040 52570 202500
rect 55570 202500 60690 202620
rect 548610 202500 549270 204960
rect 55570 202490 60730 202500
rect 55570 202470 59960 202490
rect 55550 202420 59960 202470
rect 46040 201770 52570 202040
rect 44080 201740 52570 201770
rect 44080 201560 46260 201740
rect 52270 201070 52570 201740
rect 44914 200770 44920 201070
rect 45220 200770 52570 201070
rect 52270 200130 52570 200770
rect 45014 199830 45020 200130
rect 45320 199830 52570 200130
rect 52270 199110 52570 199830
rect 56060 201090 56260 202420
rect 56590 201090 56790 202420
rect 56060 200890 56790 201090
rect 56060 199720 56260 200890
rect 57320 199720 57520 202420
rect 56060 199520 57520 199720
rect 56060 199110 56260 199520
rect 58170 199110 58370 202420
rect 545850 202320 549270 202500
rect 45444 198810 45450 199110
rect 45750 198950 52980 199110
rect 45750 198850 53000 198950
rect 45750 198810 52980 198850
rect 53170 196510 53270 198950
rect 53510 196530 53610 198880
rect 53870 196530 53970 198950
rect 53164 196410 53170 196510
rect 53270 196410 53276 196510
rect 53504 196430 53510 196530
rect 53610 196430 53616 196530
rect 53870 196424 53970 196430
rect 54230 196430 54330 198950
rect 54590 196480 54690 198950
rect 54590 196374 54690 196380
rect 54950 196430 55050 198950
rect 54230 196324 54330 196330
rect 54950 196324 55050 196330
rect 55310 196350 55410 198950
rect 56060 198910 58370 199110
rect 56060 198890 56260 198910
rect 55310 196250 55760 196350
rect 55860 196250 55866 196350
rect 18576 160310 162494 160435
rect 18576 158440 151710 160310
rect 162360 158440 162494 160310
rect 18576 158366 162494 158440
rect 171194 129980 171200 130040
rect 171260 129980 191546 130040
rect 191486 104570 191546 129980
rect 191480 104510 191486 104570
rect 191546 104510 191552 104570
rect 180444 91640 180450 91850
rect 180660 91640 181070 91850
rect 189760 91640 190905 91850
rect 191115 91640 191121 91850
rect 166148 87960 166154 88273
rect 166467 88270 181603 88273
rect 182025 88270 182075 88273
rect 183025 88270 183075 88273
rect 183604 88270 184283 88273
rect 185025 88270 185075 88273
rect 186025 88270 186075 88273
rect 187025 88270 187075 88273
rect 188025 88270 188075 88273
rect 189025 88270 189075 88273
rect 190025 88270 190075 88273
rect 166467 88150 202755 88270
rect 166467 87960 183790 88150
rect 184030 87960 202755 88150
rect 203065 87960 203071 88270
rect 181090 78165 181160 87960
rect 182090 78355 182160 87960
rect 182084 78285 182090 78355
rect 182160 78285 182166 78355
rect 183090 78245 183160 87960
rect 184090 78335 184160 87960
rect 184090 78259 184160 78265
rect 183090 78169 183160 78175
rect 179499 78095 179505 78165
rect 179575 78095 181160 78165
rect 185090 78165 185160 87960
rect 186090 78545 186160 87960
rect 187090 78655 187160 87960
rect 187090 78579 187160 78585
rect 186090 78469 186160 78475
rect 188090 78325 188160 87960
rect 189090 78495 189160 87960
rect 189090 78419 189160 78425
rect 190090 78435 190160 87960
rect 190090 78359 190160 78365
rect 188090 78249 188160 78255
rect 185090 78089 185160 78095
<< via1 >>
rect 22560 691070 26520 692780
rect 36060 687790 39510 689470
rect 26663 682328 27687 683632
rect 29716 682806 30585 683675
rect 31111 683151 31609 683649
rect 57316 224245 59385 226314
rect 44290 203870 46040 204950
rect 55880 204740 57195 204930
rect 53774 204532 53844 204538
rect 53774 204462 53780 204532
rect 53780 204462 53844 204532
rect 53774 204456 53844 204462
rect 49580 204350 49640 204410
rect 44290 203470 53490 203870
rect 44290 201770 46040 203470
rect 60690 202500 548610 204960
rect 44920 200770 45220 201070
rect 45020 199830 45320 200130
rect 45450 198810 45750 199110
rect 53170 196410 53270 196510
rect 53510 196430 53610 196530
rect 53870 196430 53970 196530
rect 54230 196330 54330 196430
rect 54590 196380 54690 196480
rect 54950 196330 55050 196430
rect 55760 196250 55860 196350
rect 151710 158440 162360 160310
rect 171200 129980 171260 130040
rect 191486 104510 191546 104570
rect 180450 91640 180660 91850
rect 190905 91640 191115 91850
rect 166154 87960 166467 88273
rect 202755 87960 203065 88270
rect 182090 78285 182160 78355
rect 184090 78265 184160 78335
rect 183090 78175 183160 78245
rect 179505 78095 179575 78165
rect 187090 78585 187160 78655
rect 186090 78475 186160 78545
rect 189090 78425 189160 78495
rect 190090 78365 190160 78435
rect 188090 78255 188160 78325
rect 185090 78095 185160 78165
<< metal2 >>
rect 165590 697195 165599 699685
rect 168089 697195 168098 699685
rect 24140 692850 26600 692870
rect 22490 692780 26600 692850
rect 22490 691070 22560 692780
rect 26520 691070 26600 692780
rect 22490 690940 26600 691070
rect 2500 690175 5000 690600
rect 24140 690410 24300 690940
rect 24830 690410 26600 690940
rect 2500 690080 25285 690175
rect 795 690030 25500 690080
rect 2500 688525 25285 690030
rect 2500 685237 5000 688525
rect 2496 682747 2505 685237
rect 4995 682747 5004 685237
rect 10250 684986 10390 684990
rect 26505 684986 26585 684990
rect 10200 684981 26590 684986
rect 10200 684901 26505 684981
rect 26585 684901 26590 684981
rect 10200 684896 26590 684901
rect 10250 683795 10390 684896
rect 26505 684892 26585 684896
rect 26750 684545 26840 689715
rect 27260 685805 27350 689705
rect 27260 685715 28325 685805
rect 14975 684455 26840 684545
rect 10246 683665 10255 683795
rect 10385 683665 10394 683795
rect 10250 683660 10390 683665
rect 2500 682742 5000 682747
rect 14975 681795 15065 684455
rect 26663 683632 27687 683641
rect 26657 682328 26663 683632
rect 27687 682328 27693 683632
rect 26663 682319 27687 682328
rect 14975 681670 15065 681705
rect 5720 681055 6040 681100
rect 28235 681055 28325 685715
rect 29716 683675 30585 683684
rect 29710 682806 29716 683675
rect 30585 682806 30591 683675
rect 31111 683649 31609 683658
rect 31105 683151 31111 683649
rect 31609 683151 31615 683649
rect 31111 683142 31609 683151
rect 29716 682797 30585 682806
rect 5195 680965 28325 681055
rect 5720 678115 6040 680965
rect 14975 680400 15065 680450
rect 14971 680320 14980 680400
rect 15060 680320 15069 680400
rect 5716 677805 5725 678115
rect 6035 677805 6044 678115
rect 5720 677800 6040 677805
rect 14975 672355 15065 680320
rect 14966 672265 14975 672355
rect 15065 672265 15074 672355
rect 32590 206138 32670 689740
rect 33290 207748 33370 689730
rect 33290 207692 33302 207748
rect 33358 207692 33370 207748
rect 33290 207480 33370 207692
rect 32590 206082 32592 206138
rect 32648 206082 32670 206138
rect 32590 193540 32670 206082
rect 34420 199300 34500 689730
rect 35960 689470 39580 689550
rect 35960 687790 36060 689470
rect 39510 689460 39580 689470
rect 39510 689345 42700 689460
rect 39510 687790 40195 689345
rect 35960 687690 40195 687790
rect 35990 686895 40195 687690
rect 42645 686900 42700 689345
rect 42645 686895 42650 686900
rect 35990 686890 42650 686895
rect 40195 686886 42645 686890
rect 40343 339375 40352 339445
rect 40422 339375 49997 339445
rect 44080 204950 46260 205280
rect 44080 201770 44290 204950
rect 46040 204150 46260 204950
rect 49927 204532 49997 339375
rect 57316 226314 59385 226320
rect 57312 224250 57316 226309
rect 59385 224250 59389 226309
rect 57316 224239 59385 224245
rect 54101 211840 54110 211900
rect 54170 211840 54179 211900
rect 54120 204770 54160 211840
rect 54500 209860 54509 209920
rect 54569 209860 54578 209920
rect 54519 204770 54559 209860
rect 54935 207480 54944 207540
rect 55004 207480 55013 207540
rect 54954 204770 54994 207480
rect 56530 205690 56590 205699
rect 56530 205621 56590 205630
rect 55389 205100 55429 205110
rect 56540 205100 56580 205621
rect 55389 205060 56590 205100
rect 55389 204620 55429 205060
rect 545850 205030 549270 205460
rect 60625 204980 549270 205030
rect 55830 204960 549270 204980
rect 55830 204930 60690 204960
rect 55830 204740 55880 204930
rect 60615 204740 60690 204930
rect 55830 204710 60690 204740
rect 53774 204538 53844 204544
rect 49927 204462 53774 204532
rect 53774 204450 53844 204456
rect 49580 204410 49640 204419
rect 49574 204350 49580 204410
rect 49640 204350 49646 204410
rect 49580 204341 49640 204350
rect 46040 203890 53610 204150
rect 46040 203870 53620 203890
rect 53490 203470 53620 203870
rect 46040 203410 53620 203470
rect 46040 201770 46260 203410
rect 53160 203085 53200 203090
rect 53160 203055 53949 203085
rect 53160 202790 53200 203055
rect 54350 203000 54390 203090
rect 55224 203082 55254 203085
rect 54789 203055 54819 203080
rect 53500 202998 53560 203000
rect 53493 202942 53502 202998
rect 53558 202942 53567 202998
rect 53840 202960 54390 203000
rect 54625 203025 54819 203055
rect 53500 202760 53560 202942
rect 53840 202790 53880 202960
rect 54231 202860 54287 202867
rect 54170 202858 54300 202860
rect 54170 202802 54231 202858
rect 54287 202802 54300 202858
rect 54625 202830 54655 203025
rect 54840 202968 54900 202970
rect 54833 202912 54842 202968
rect 54898 202912 54907 202968
rect 54170 202730 54300 202802
rect 54520 202790 54655 202830
rect 54525 202785 54655 202790
rect 54840 202770 54900 202912
rect 55208 202785 55254 203082
rect 55530 202948 55590 202950
rect 55523 202892 55532 202948
rect 55588 202892 55597 202948
rect 55530 202770 55590 202892
rect 60625 202500 60690 204710
rect 548610 202500 549270 204960
rect 545850 202320 549270 202500
rect 44080 201560 46260 201770
rect 44920 201070 45220 201076
rect 44911 200770 44920 201070
rect 45220 200770 45229 201070
rect 44920 200764 45220 200770
rect 45020 200130 45320 200136
rect 45011 199830 45020 200130
rect 45320 199830 45329 200130
rect 45020 199824 45320 199830
rect 48460 199310 51040 199330
rect 48460 199300 48480 199310
rect 34420 199220 48480 199300
rect 34420 124690 34500 199220
rect 48460 199180 48480 199220
rect 51020 199180 51040 199310
rect 48460 199170 51040 199180
rect 45450 199110 45750 199116
rect 45441 198810 45450 199110
rect 45750 198810 45759 199110
rect 45450 198804 45750 198810
rect 53510 196530 53610 196536
rect 53870 196530 53970 196539
rect 53170 196510 53270 196516
rect 53161 196410 53170 196510
rect 53270 196410 53279 196510
rect 53501 196430 53510 196530
rect 53610 196430 53619 196530
rect 53864 196430 53870 196530
rect 53970 196430 53976 196530
rect 54590 196480 54690 196489
rect 54584 196470 54590 196480
rect 54200 196430 54350 196460
rect 53510 196424 53610 196430
rect 53870 196421 53970 196430
rect 53170 196404 53270 196410
rect 54200 196330 54230 196430
rect 54330 196330 54350 196430
rect 54581 196380 54590 196470
rect 54690 196470 54696 196480
rect 54690 196380 54699 196470
rect 54950 196430 55050 196439
rect 54590 196371 54690 196380
rect 54944 196330 54950 196430
rect 55050 196330 55056 196430
rect 55760 196350 55860 196356
rect 54200 196280 54350 196330
rect 54950 196321 55050 196330
rect 55751 196250 55760 196350
rect 55860 196250 55869 196350
rect 55760 196244 55860 196250
rect 151670 160310 162410 160340
rect 151670 158440 151710 160310
rect 162360 158440 162410 160310
rect 151670 158410 162410 158440
rect 184216 153583 184225 153700
rect 184342 153583 184351 153700
rect 180381 152314 180536 152323
rect 180381 152150 180536 152159
rect 171200 130040 171260 130046
rect 171191 129980 171200 130040
rect 171260 129980 171269 130040
rect 171200 129974 171260 129980
rect 34190 124590 34820 124690
rect 34190 119850 34290 124590
rect 34180 119700 34290 119850
rect 34680 119700 34820 124590
rect 34180 119290 34820 119700
rect 180428 116224 180488 152150
rect 182353 145677 182487 145686
rect 182353 145534 182487 145543
rect 180428 116164 182360 116224
rect 4150 115910 178656 116050
rect 4150 81661 4290 115910
rect 178516 101670 178656 115910
rect 182300 104038 182360 116164
rect 182293 103982 182302 104038
rect 182358 103982 182367 104038
rect 182300 103980 182360 103982
rect 182400 102733 182440 145534
rect 182684 141210 182847 141219
rect 182684 141038 182847 141047
rect 182735 104274 182795 141038
rect 182948 135992 183145 136001
rect 182948 135786 183145 135795
rect 182728 104218 182737 104274
rect 182793 104218 182802 104274
rect 182735 104216 182795 104218
rect 183026 102989 183066 135786
rect 184253 130386 184313 153583
rect 192704 152350 192871 152359
rect 192704 152174 192871 152183
rect 185361 146684 185480 146693
rect 185361 145768 185480 146565
rect 184253 130326 185360 130386
rect 183122 127739 183279 127748
rect 183122 125375 183279 127582
rect 183170 103962 183230 125375
rect 183353 123800 183461 123809
rect 183353 123683 183461 123692
rect 183163 103906 183172 103962
rect 183228 103906 183237 103962
rect 183170 103904 183230 103906
rect 182835 102949 183066 102989
rect 182835 102705 182875 102949
rect 183387 102783 183427 123683
rect 183569 120059 183701 120278
rect 183569 119161 183701 119927
rect 183605 104150 183665 119161
rect 184250 117486 184370 117495
rect 184250 117191 184370 117366
rect 184290 106769 184330 117191
rect 183705 106729 184330 106769
rect 183602 104008 183668 104150
rect 183598 103952 183672 104008
rect 183602 103587 183668 103952
rect 183598 103531 183607 103587
rect 183663 103531 183672 103587
rect 183602 103526 183668 103531
rect 183270 102743 183427 102783
rect 183705 102698 183745 106729
rect 185300 103639 185360 130326
rect 185293 103583 185302 103639
rect 185358 103583 185367 103639
rect 185300 103581 185360 103583
rect 185400 102714 185440 145768
rect 185941 141836 186059 141845
rect 185941 141303 186059 141718
rect 185970 104892 186030 141303
rect 186811 136373 186871 136382
rect 186811 136304 186871 136313
rect 185735 104890 186030 104892
rect 185728 104834 185737 104890
rect 185793 104834 186030 104890
rect 185735 104832 186030 104834
rect 186821 104421 186861 136304
rect 187094 128327 187196 128336
rect 187094 127496 187196 128225
rect 185835 104381 186861 104421
rect 185835 102708 185875 104381
rect 186432 104199 186488 104206
rect 187115 104199 187175 127496
rect 187326 123736 187409 123745
rect 187326 123644 187409 123653
rect 186430 104197 187175 104199
rect 186430 104141 186432 104197
rect 186488 104141 187175 104197
rect 186430 104139 187175 104141
rect 186432 104132 186488 104139
rect 187347 104067 187387 123644
rect 187567 120881 187673 120890
rect 187567 120766 187673 120775
rect 186270 104027 187387 104067
rect 186270 102740 186310 104027
rect 186590 103802 186680 103806
rect 186585 103797 187539 103802
rect 186585 103707 186590 103797
rect 186680 103785 187539 103797
rect 187587 103785 187653 120766
rect 187976 117391 188036 117400
rect 187976 117322 188036 117331
rect 186680 103719 187653 103785
rect 186680 103707 187539 103719
rect 186585 103702 187539 103707
rect 186590 103698 186680 103702
rect 187986 103366 188026 117322
rect 192757 105059 192817 152174
rect 195086 146728 195188 146737
rect 195086 145974 195188 146626
rect 188300 104999 192817 105059
rect 188300 103698 188360 104999
rect 195117 104934 195157 145974
rect 197541 141810 197550 141870
rect 197610 141810 197619 141870
rect 188400 104894 195157 104934
rect 188293 103642 188302 103698
rect 188358 103642 188367 103698
rect 188300 103640 188360 103642
rect 186705 103326 188026 103366
rect 186705 102724 186745 103326
rect 188400 102699 188440 104894
rect 192842 104760 192898 104767
rect 197550 104760 197610 141810
rect 201061 136700 201070 136760
rect 201130 136700 201139 136760
rect 192840 104758 197610 104760
rect 192840 104702 192842 104758
rect 192898 104702 197610 104758
rect 192840 104700 197610 104702
rect 192842 104693 192898 104700
rect 191486 104570 191546 104576
rect 191479 104512 191486 104568
rect 191546 104512 191553 104568
rect 191486 104504 191546 104510
rect 201080 104450 201120 136700
rect 188835 104410 201120 104450
rect 205240 128370 205300 128379
rect 188835 102650 188875 104410
rect 189172 104130 189228 104137
rect 205240 104130 205300 128310
rect 206310 124450 206370 124459
rect 206310 124381 206370 124390
rect 189170 104128 205300 104130
rect 189170 104072 189172 104128
rect 189228 104072 205300 104128
rect 189170 104070 205300 104072
rect 189172 104063 189228 104070
rect 206320 103400 206360 124381
rect 189270 103360 206360 103400
rect 208020 120760 208080 120769
rect 189270 102720 189310 103360
rect 189607 103140 189663 103147
rect 208020 103140 208080 120700
rect 212530 105820 212590 105829
rect 212530 105751 212590 105760
rect 189605 103138 208080 103140
rect 189605 103082 189607 103138
rect 189663 103082 208080 103138
rect 189605 103080 208080 103082
rect 189607 103073 189663 103080
rect 212540 102757 212580 105751
rect 189705 102717 212580 102757
rect 10250 92690 10390 92699
rect 10390 92550 178146 92690
rect 10250 92541 10390 92550
rect 10954 91069 11066 91076
rect 179908 91069 180045 92316
rect 180450 91850 180660 91856
rect 190905 91850 191115 91856
rect 180441 91640 180450 91850
rect 180660 91640 180669 91850
rect 190896 91640 190905 91850
rect 191115 91640 191124 91850
rect 180450 91634 180660 91640
rect 190905 91634 191115 91640
rect 10930 90932 180045 91069
rect 4150 81559 4179 81661
rect 4281 81559 4290 81661
rect 4150 81460 4290 81559
rect 10954 39756 11066 90932
rect 166154 88273 166467 88279
rect 166145 87960 166154 88273
rect 166467 87960 166476 88273
rect 166154 87954 166467 87960
rect 184215 80148 184275 80150
rect 187215 80148 187275 80150
rect 184208 80092 184217 80148
rect 184273 80092 184282 80148
rect 187208 80092 187217 80148
rect 187273 80092 187282 80148
rect 182915 79978 182975 79980
rect 182908 79922 182917 79978
rect 182973 79922 182982 79978
rect 181895 79778 181955 79780
rect 181888 79722 181897 79778
rect 181953 79722 181962 79778
rect 179505 78165 179575 78171
rect 179496 78095 179505 78165
rect 179575 78095 179584 78165
rect 179505 78089 179575 78095
rect 1774 39644 11066 39756
rect 1774 38439 1886 39644
rect 1774 38337 1779 38439
rect 1881 38337 1886 38439
rect 1774 38332 1886 38337
rect 1779 38328 1881 38332
rect 157721 29354 157730 29466
rect 157842 29354 157851 29466
rect 75730 26498 75790 26500
rect 75723 26442 75732 26498
rect 75788 26442 75797 26498
rect 75730 10626 75790 26442
rect 72344 10514 155478 10626
rect 75730 10320 75790 10514
rect 69764 8646 69876 8655
rect 68454 8534 69764 8646
rect 69876 8534 151932 8646
rect 69764 8525 69876 8534
rect 66364 7086 66476 7095
rect 64844 6974 66364 7086
rect 66476 6974 148386 7086
rect 66364 6965 66476 6974
rect 62874 5706 62986 5715
rect 56514 5594 62874 5706
rect 62986 5594 144840 5706
rect 62874 5585 62986 5594
rect 55244 4376 55356 4385
rect 54284 4264 55244 4376
rect 55356 4264 141294 4376
rect 55244 4255 55356 4264
rect 52334 3346 52446 3355
rect 50394 3234 52334 3346
rect 52446 3234 137748 3346
rect 52334 3225 52446 3234
rect 49534 2266 49646 2275
rect 47484 2154 49534 2266
rect 49646 2154 134202 2266
rect 49534 2145 49646 2154
rect 46414 1726 46526 1735
rect 44074 1614 46414 1726
rect 46526 1614 130656 1726
rect 46414 1605 46526 1614
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 1614
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 2154
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 3234
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 4264
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 5594
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 6974
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 8534
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 10514
rect 156548 -800 156660 480
rect 157730 -800 157842 29354
rect 161276 28706 161388 28715
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 28594
rect 181895 28280 181955 79722
rect 182235 79688 182295 79690
rect 182228 79632 182237 79688
rect 182293 79632 182302 79688
rect 182090 78355 182160 78361
rect 182081 78285 182090 78355
rect 182160 78285 182169 78355
rect 182090 78279 182160 78285
rect 164830 28256 181955 28280
rect 164822 28220 181955 28256
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 28220
rect 168368 27630 168480 27816
rect 182235 27630 182295 79632
rect 168368 27570 182295 27630
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 27570
rect 171914 27080 172026 27096
rect 182577 27080 182633 27087
rect 171860 27078 182635 27080
rect 171860 27022 182577 27078
rect 182633 27022 182635 27078
rect 171860 27020 182635 27022
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 27020
rect 182577 27013 182633 27020
rect 175460 26320 175572 26336
rect 182915 26320 182975 79922
rect 183255 79568 183315 79570
rect 183248 79512 183257 79568
rect 183313 79512 183322 79568
rect 183090 78245 183160 78254
rect 183084 78175 183090 78245
rect 183160 78175 183166 78245
rect 183090 78166 183160 78175
rect 175410 26260 182975 26320
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 26260
rect 179006 25400 179118 25416
rect 183255 25400 183315 79512
rect 184090 78335 184160 78344
rect 184084 78265 184090 78335
rect 184160 78265 184166 78335
rect 184090 78256 184160 78265
rect 178830 25340 183315 25400
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 25340
rect 182552 23676 182664 23685
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 23564
rect 184215 1496 184275 80092
rect 185915 79978 185975 79980
rect 185908 79922 185917 79978
rect 185973 79922 185982 79978
rect 184895 79778 184955 79780
rect 184888 79722 184897 79778
rect 184953 79722 184962 79778
rect 184895 3170 184955 79722
rect 185235 79688 185295 79690
rect 185228 79632 185237 79688
rect 185293 79632 185302 79688
rect 185090 78165 185160 78174
rect 185084 78095 185090 78165
rect 185160 78095 185166 78165
rect 185090 78086 185160 78095
rect 185235 3690 185295 79632
rect 185915 4900 185975 79922
rect 186255 79568 186315 79570
rect 186248 79512 186257 79568
rect 186313 79512 186322 79568
rect 186090 78545 186160 78554
rect 186084 78475 186090 78545
rect 186160 78475 186166 78545
rect 186090 78466 186160 78475
rect 186255 5760 186315 79512
rect 187090 78655 187160 78664
rect 187084 78585 187090 78655
rect 187160 78585 187166 78655
rect 187090 78576 187160 78585
rect 187215 7050 187275 80092
rect 188915 79978 188975 79980
rect 188908 79922 188917 79978
rect 188973 79922 188982 79978
rect 187895 79778 187955 79780
rect 187888 79722 187897 79778
rect 187953 79722 187962 79778
rect 187895 7790 187955 79722
rect 188235 79688 188295 79690
rect 188228 79632 188237 79688
rect 188293 79632 188302 79688
rect 188090 78325 188160 78334
rect 188084 78255 188090 78325
rect 188160 78255 188166 78325
rect 188090 78246 188160 78255
rect 188235 8640 188295 79632
rect 188915 9140 188975 79922
rect 189255 79568 189315 79570
rect 189248 79512 189257 79568
rect 189313 79512 189322 79568
rect 189090 78495 189160 78504
rect 189084 78425 189090 78495
rect 189160 78425 189166 78495
rect 189090 78416 189160 78425
rect 189255 9410 189315 79512
rect 190090 78435 190160 78444
rect 190084 78365 190090 78435
rect 190160 78365 190166 78435
rect 190090 78356 190160 78365
rect 191205 73062 191368 92217
rect 202755 88270 203065 88276
rect 202746 87960 202755 88270
rect 203065 87960 203074 88270
rect 202755 87954 203065 87960
rect 191205 72899 549680 73062
rect 239279 9694 239288 9806
rect 239400 9694 239409 9806
rect 235742 9410 235854 9486
rect 189255 9350 236220 9410
rect 188915 9080 233210 9140
rect 188577 8940 188633 8947
rect 228650 8940 228762 9030
rect 188575 8938 228762 8940
rect 188575 8882 188577 8938
rect 188633 8882 228762 8938
rect 188575 8880 228762 8882
rect 188577 8873 188633 8880
rect 225104 8640 225216 8696
rect 188235 8580 226120 8640
rect 221558 7790 221670 7796
rect 187895 7730 222040 7790
rect 218012 7286 218124 7295
rect 218003 7184 218012 7286
rect 218124 7184 218133 7286
rect 214466 7050 214578 7086
rect 187215 6990 215300 7050
rect 210920 6358 211032 6486
rect 210920 6302 210962 6358
rect 211018 6302 211032 6358
rect 207374 5760 207486 5776
rect 186255 5700 208070 5760
rect 203194 4900 203940 4916
rect 185915 4840 203940 4900
rect 203194 4804 203940 4840
rect 185577 4450 185633 4457
rect 185575 4448 200510 4450
rect 185575 4392 185577 4448
rect 185633 4392 200510 4448
rect 185575 4390 200510 4392
rect 185577 4383 185633 4390
rect 196736 3690 196848 3756
rect 185235 3630 196848 3690
rect 193190 3170 193302 3186
rect 184895 3110 193302 3170
rect 184557 2500 184613 2507
rect 189644 2500 189756 2516
rect 184555 2498 189756 2500
rect 184555 2442 184557 2498
rect 184613 2442 189756 2498
rect 184555 2440 189756 2442
rect 184557 2433 184613 2440
rect 184215 1384 186210 1496
rect 184215 1280 184275 1384
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 1384
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 2440
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 3110
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 3630
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 4390
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 4804
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 5700
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 6302
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 6990
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 7174
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 7730
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 8580
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 8880
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 9080
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 9350
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 9694
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 72899
rect 551336 10576 551448 10936
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 10464
rect 576158 9736 576270 10116
rect 576149 9624 576158 9736
rect 576270 9624 576279 9736
rect 558428 7876 558540 8316
rect 554882 6156 554994 7226
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 6044
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 7764
rect 572612 6556 572724 6686
rect 561974 6076 562086 6356
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 5964
rect 565520 6306 565632 6406
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 6194
rect 569066 6286 569178 6466
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 6174
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 6444
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 9624
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 165599 697195 168089 699685
rect 22560 691070 26520 692780
rect 24300 690410 24830 690940
rect 2505 682747 4995 685237
rect 26505 684901 26585 684981
rect 10255 683665 10385 683795
rect 26663 682328 27687 683632
rect 14975 681705 15065 681795
rect 29716 682806 30585 683675
rect 31111 683151 31609 683649
rect 14980 680320 15060 680400
rect 5725 677805 6035 678115
rect 14975 672265 15065 672355
rect 33302 207692 33358 207748
rect 32592 206082 32648 206138
rect 40195 686895 42645 689345
rect 40352 339375 40422 339445
rect 44290 203870 46040 204950
rect 57321 224250 59380 226309
rect 54110 211840 54170 211900
rect 54509 209860 54569 209920
rect 54944 207480 55004 207540
rect 56530 205630 56590 205690
rect 55880 204740 57195 204930
rect 57195 204740 60615 204930
rect 49580 204350 49640 204410
rect 44290 203470 53490 203870
rect 44290 201770 46040 203470
rect 53502 202942 53558 202998
rect 54231 202802 54287 202858
rect 54842 202912 54898 202968
rect 55532 202892 55588 202948
rect 60690 202500 548610 204960
rect 44920 200770 45220 201070
rect 45020 199830 45320 200130
rect 48480 199180 51020 199310
rect 45450 198810 45750 199110
rect 53170 196410 53270 196510
rect 53510 196430 53610 196530
rect 53870 196430 53970 196530
rect 54230 196330 54330 196430
rect 54590 196380 54690 196480
rect 54950 196330 55050 196430
rect 55760 196250 55860 196350
rect 151710 158440 162360 160310
rect 184225 153583 184342 153700
rect 180381 152159 180536 152314
rect 171200 129980 171260 130040
rect 34290 119700 34680 124590
rect 182353 145543 182487 145677
rect 182302 103982 182358 104038
rect 182684 141047 182847 141210
rect 182948 135795 183145 135992
rect 182737 104218 182793 104274
rect 192704 152183 192871 152350
rect 185361 146565 185480 146684
rect 183122 127582 183279 127739
rect 183353 123692 183461 123800
rect 183172 103906 183228 103962
rect 183569 119927 183701 120059
rect 184250 117366 184370 117486
rect 183607 103531 183663 103587
rect 185302 103583 185358 103639
rect 185941 141718 186059 141836
rect 186811 136313 186871 136373
rect 185737 104834 185793 104890
rect 187094 128225 187196 128327
rect 187326 123653 187409 123736
rect 186432 104141 186488 104197
rect 187567 120775 187673 120881
rect 186590 103707 186680 103797
rect 187976 117331 188036 117391
rect 195086 146626 195188 146728
rect 197550 141810 197610 141870
rect 188302 103642 188358 103698
rect 201070 136700 201130 136760
rect 192842 104702 192898 104758
rect 191488 104512 191544 104568
rect 205240 128310 205300 128370
rect 206310 124390 206370 124450
rect 189172 104072 189228 104128
rect 208020 120700 208080 120760
rect 212530 105760 212590 105820
rect 189607 103082 189663 103138
rect 10250 92550 10390 92690
rect 180450 91640 180660 91850
rect 190905 91640 191115 91850
rect 4179 81559 4281 81661
rect 166154 87960 166467 88273
rect 184217 80092 184273 80148
rect 187217 80092 187273 80148
rect 182917 79922 182973 79978
rect 181897 79722 181953 79778
rect 179505 78095 179575 78165
rect 1779 38337 1881 38439
rect 157730 29354 157842 29466
rect 75732 26442 75788 26498
rect 69764 8534 69876 8646
rect 66364 6974 66476 7086
rect 62874 5594 62986 5706
rect 55244 4264 55356 4376
rect 52334 3234 52446 3346
rect 49534 2154 49646 2266
rect 46414 1614 46526 1726
rect 161276 28594 161388 28706
rect 182237 79632 182293 79688
rect 182090 78285 182160 78355
rect 182577 27022 182633 27078
rect 183257 79512 183313 79568
rect 183090 78175 183160 78245
rect 184090 78265 184160 78335
rect 182552 23564 182664 23676
rect 185917 79922 185973 79978
rect 184897 79722 184953 79778
rect 185237 79632 185293 79688
rect 185090 78095 185160 78165
rect 186257 79512 186313 79568
rect 186090 78475 186160 78545
rect 187090 78585 187160 78655
rect 188917 79922 188973 79978
rect 187897 79722 187953 79778
rect 188237 79632 188293 79688
rect 188090 78255 188160 78325
rect 189257 79512 189313 79568
rect 189090 78425 189160 78495
rect 190090 78365 190160 78435
rect 202755 87960 203065 88270
rect 239288 9694 239400 9806
rect 188577 8882 188633 8938
rect 218012 7174 218124 7286
rect 210962 6302 211018 6358
rect 185577 4392 185633 4448
rect 184557 2442 184613 2498
rect 551336 10464 551448 10576
rect 576158 9624 576270 9736
rect 558428 7764 558540 7876
rect 554882 6044 554994 6156
rect 561974 5964 562086 6076
rect 565520 6194 565632 6306
rect 569066 6174 569178 6286
rect 572612 6444 572724 6556
<< metal3 >>
rect 16194 703310 21194 704800
rect 16194 702300 27065 703310
rect 18694 701630 27065 702300
rect 68194 702300 73194 704800
rect 120194 702740 125194 704800
rect 75620 702300 125194 702740
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702310 470394 704800
rect 420980 702300 470394 702310
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 68194 701860 70694 702300
rect 18694 699900 27220 701630
rect 68140 700540 70694 701860
rect 29770 699960 70694 700540
rect 24590 695880 25050 695886
rect 22584 695320 22590 695780
rect 23050 695320 23056 695780
rect 23590 695770 24050 695776
rect 22590 692850 23050 695320
rect 23590 692850 24050 695310
rect 24590 692870 25050 695420
rect 25590 695880 26050 695886
rect 25590 692870 26050 695420
rect 24140 692850 26600 692870
rect 22490 692780 26600 692850
rect 22490 691070 22560 692780
rect 26520 691070 26600 692780
rect 22490 690940 26600 691070
rect 22490 690410 24300 690940
rect 24830 690410 26600 690940
rect 27020 690560 27220 699900
rect 27530 699760 70694 699960
rect 27530 690590 27730 699760
rect 29770 699360 70694 699760
rect 75620 701700 124910 702300
rect 29770 699320 70270 699360
rect 75620 698120 76660 701700
rect 319171 701179 321669 701185
rect 164800 700260 168840 700320
rect 28410 697080 76660 698120
rect 77320 699689 168890 700260
rect 218481 700130 220979 700135
rect 77320 699240 165595 699689
rect -800 685237 5000 685242
rect -800 682747 2505 685237
rect 4995 682747 5000 685237
rect 10250 683799 10390 683800
rect 10245 683661 10251 683799
rect 10389 683661 10395 683799
rect 10250 683660 10390 683661
rect -800 682742 5000 682747
rect -800 680242 1700 682742
rect 14970 681795 15070 681800
rect 14970 681705 14975 681795
rect 15065 681705 15070 681795
rect 14970 681700 15070 681705
rect 14975 680400 15065 681700
rect 14975 680320 14980 680400
rect 15060 680320 15065 680400
rect 14975 680315 15065 680320
rect 22490 680270 24950 690410
rect 28410 690390 29450 697080
rect 77320 695140 78340 699240
rect 164800 697400 165595 699240
rect 165589 697191 165595 697400
rect 168093 699240 168890 699689
rect 215230 700129 220980 700130
rect 215230 699305 218481 700129
rect 168093 697400 168840 699240
rect 172955 698835 218481 699305
rect 168093 697191 168099 697400
rect 165594 697190 168094 697191
rect 30220 694120 78340 695140
rect 30220 690370 31240 694120
rect 172955 693615 173425 698835
rect 215230 697631 218481 698835
rect 220979 697631 220980 700129
rect 215230 697630 220980 697631
rect 224425 699655 319171 700125
rect 218481 697625 220979 697630
rect 32150 693145 173425 693615
rect 32150 691050 32620 693145
rect 33300 692645 33770 692675
rect 224425 692645 224895 699655
rect 319171 698675 321669 698681
rect 33300 692175 224895 692645
rect 33300 691000 33770 692175
rect 34660 691430 35130 691620
rect 415560 691430 418060 702300
rect 34660 690960 418060 691430
rect 415560 690760 418060 690960
rect 420980 699810 467894 702300
rect 26500 684981 26590 689773
rect 26500 684901 26505 684981
rect 26585 684901 26590 684981
rect 26500 684896 26590 684901
rect 29711 683675 30590 683680
rect 29711 683670 29716 683675
rect 30585 683670 30590 683675
rect 26658 683632 27692 683637
rect 26658 683627 26663 683632
rect 27687 683627 27692 683632
rect 31106 683649 31614 683654
rect 31106 683644 31111 683649
rect 31609 683644 31614 683649
rect 31106 683140 31614 683146
rect 29711 682795 30590 682801
rect 26658 682317 27692 682323
rect 22484 678880 22490 680270
rect 5720 678115 6040 678120
rect 5720 677805 5725 678115
rect 6035 677805 6040 678115
rect 5720 673659 6040 677805
rect 18410 677810 22490 678880
rect 24950 677810 24956 680270
rect 18410 676420 24950 677810
rect 5715 673341 5721 673659
rect 6039 673341 6045 673659
rect 5720 673340 6040 673341
rect 14970 672355 14980 672360
rect 14970 672265 14975 672355
rect 14970 672260 14980 672265
rect 15070 672260 15076 672360
rect 18410 648642 20870 676420
rect -800 646182 20870 648642
rect -800 643842 1660 646182
rect -800 637210 1660 638642
rect -800 634750 19000 637210
rect 21460 634750 21466 637210
rect -800 633842 1660 634750
rect -800 562060 1660 564242
rect -800 559600 14060 562060
rect 16520 559600 16526 562060
rect -800 559442 1660 559600
rect -800 552210 1660 554242
rect -800 549750 14400 552210
rect 16860 549750 16866 552210
rect -800 549442 1660 549750
rect 35680 511660 35880 690760
rect 36240 689349 42840 689740
rect 36240 686891 40191 689349
rect 42649 686891 42840 689349
rect 420980 686930 423480 699810
rect 510594 698400 513054 702340
rect 566594 702300 571594 704800
rect 569270 699299 569590 702300
rect 569265 698981 569271 699299
rect 569589 698981 569595 699299
rect 569270 698980 569590 698981
rect 36240 686560 42840 686891
rect 1360 511642 35880 511660
rect -800 511530 35880 511642
rect 1360 511460 35880 511530
rect 35680 510910 35880 511460
rect 46460 684430 423480 686930
rect 426710 695940 513054 698400
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 40347 339445 40427 339450
rect 10035 339375 40352 339445
rect 40422 339375 40427 339445
rect 10375 338754 10487 339375
rect 40347 339370 40427 339375
rect -800 338642 10552 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect -800 295420 36783 295532
rect 36895 295420 36901 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect -800 252398 30075 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect 29941 250039 30053 252398
rect 29941 249971 29956 250039
rect 30024 249971 30053 250039
rect 29941 249942 30053 249971
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect -800 214888 1660 219688
rect 46460 215520 48960 684430
rect 426710 679010 429170 695940
rect 404020 678815 429170 679010
rect 57316 676746 429170 678815
rect 582300 677984 584800 682984
rect 57316 226309 59385 676746
rect 404020 676550 429170 676746
rect 576090 644330 584800 644584
rect 576030 639784 584800 644330
rect 576030 634584 580530 639784
rect 576030 632260 584800 634584
rect 57316 224250 57321 226309
rect 59380 224250 59385 226309
rect 57316 223050 59385 224250
rect 546150 629800 584800 632260
rect 46460 213020 52500 215520
rect -800 204888 1660 209688
rect 33297 207750 33363 207753
rect 33297 207748 50340 207750
rect 33297 207692 33302 207748
rect 33358 207692 50340 207748
rect 33297 207690 50340 207692
rect 33297 207687 33363 207690
rect 32550 206142 32700 206170
rect 32550 206078 32588 206142
rect 32652 206078 32700 206142
rect 32550 206040 32700 206078
rect 43890 204950 46350 205720
rect 43890 204858 44290 204950
rect 24944 203217 24950 204858
rect 26591 203217 44290 204858
rect 46040 204150 46350 204950
rect 49500 204415 49710 204500
rect 49500 204351 49575 204415
rect 49645 204351 49710 204415
rect 50280 204460 50340 207690
rect 51420 204630 51480 213020
rect 54050 211905 54210 211940
rect 54050 211900 54111 211905
rect 54050 211840 54110 211900
rect 54050 211835 54111 211840
rect 54175 211835 54210 211905
rect 54050 211760 54210 211835
rect 54480 209925 54640 209970
rect 54480 209920 54510 209925
rect 54480 209860 54509 209920
rect 54480 209855 54510 209860
rect 54574 209855 54640 209925
rect 54480 209840 54640 209855
rect 54870 207545 55100 207570
rect 54870 207540 54945 207545
rect 54870 207480 54944 207540
rect 54870 207475 54945 207480
rect 55009 207475 55100 207545
rect 54870 207390 55100 207475
rect 546150 206970 548610 629800
rect 582340 629784 584800 629800
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583280 313652 584800 313764
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect 56480 205695 56640 205750
rect 56480 205631 56525 205695
rect 56595 205631 56640 205695
rect 56480 205630 56530 205631
rect 56590 205630 56640 205631
rect 56480 205590 56640 205630
rect 546150 205030 549530 206970
rect 60625 204970 549530 205030
rect 53760 204960 549530 204970
rect 53760 204930 60690 204960
rect 53760 204820 55880 204930
rect 53670 204740 55880 204820
rect 60615 204740 60690 204930
rect 53670 204710 60690 204740
rect 53670 204700 55480 204710
rect 51360 204570 55530 204630
rect 50280 204400 55610 204460
rect 49500 204350 49580 204351
rect 49640 204350 49710 204351
rect 49500 204310 49710 204350
rect 46040 203890 53610 204150
rect 46040 203870 53620 203890
rect 53490 203470 53620 203870
rect 43890 201770 44290 203217
rect 46040 203410 53620 203470
rect 46040 201770 46350 203410
rect 51754 203210 53660 203270
rect 51754 203032 51814 203210
rect 51752 203026 51816 203032
rect 51752 202956 51816 202962
rect 53480 203002 53600 203020
rect 53480 202938 53498 203002
rect 53562 202938 53600 203002
rect 53480 202920 53600 202938
rect 54820 202972 54910 202990
rect 54820 202908 54838 202972
rect 54902 202908 54910 202972
rect 54820 202880 54910 202908
rect 55510 202952 55630 202990
rect 55510 202888 55528 202952
rect 55592 202888 55630 202952
rect 55510 202880 55630 202888
rect 54227 202863 54291 202868
rect 54226 202862 54292 202863
rect 54226 202860 54227 202862
rect 54170 202798 54227 202860
rect 54291 202860 54292 202862
rect 54291 202798 54300 202860
rect 54170 202730 54300 202798
rect 60625 202500 60690 204710
rect 548610 202500 549530 204960
rect 43890 201075 46350 201770
rect 59565 201630 549530 202500
rect 547970 201620 549530 201630
rect 24649 200765 25772 200771
rect 43890 200765 44915 201075
rect 45215 201070 46350 201075
rect 45220 200770 46350 201070
rect 45215 200765 46350 200770
rect 24643 199640 24649 200765
rect 25774 200135 46350 200765
rect 25774 199825 45015 200135
rect 45315 200130 46350 200135
rect 45320 199830 46350 200130
rect 45315 199825 46350 199830
rect 25774 199640 46350 199825
rect 24649 199634 25772 199640
rect 43890 199115 46350 199640
rect 49178 199490 49184 199560
rect 49254 199490 52935 199560
rect 48460 199310 51040 199330
rect 48460 199180 48480 199310
rect 51020 199240 51040 199310
rect 51020 199180 52930 199240
rect 48460 199170 51040 199180
rect 43890 198805 45445 199115
rect 45745 199110 46350 199115
rect 45750 198810 46350 199110
rect 45745 198805 46350 198810
rect 24781 197784 27239 197790
rect 43890 197784 46350 198805
rect 24775 195324 24781 197784
rect 27241 196650 46350 197784
rect 27241 196530 57890 196650
rect 27241 196510 53510 196530
rect 27241 196410 53170 196510
rect 53270 196430 53510 196510
rect 53610 196430 53870 196530
rect 53970 196480 57890 196530
rect 53970 196430 54590 196480
rect 53270 196410 54230 196430
rect 27241 196330 54230 196410
rect 54330 196380 54590 196430
rect 54690 196430 57890 196480
rect 54690 196380 54950 196430
rect 54330 196330 54950 196380
rect 55050 196355 57890 196430
rect 55050 196350 55765 196355
rect 55050 196330 55760 196350
rect 27241 196250 55760 196330
rect 27241 196245 55765 196250
rect 55865 196245 57890 196355
rect 27241 195324 57890 196245
rect 24781 195318 27239 195324
rect 43890 194190 57890 195324
rect 24930 191312 27388 191318
rect 43890 191312 46350 194190
rect 582340 191430 584800 196230
rect 24924 188852 24930 191312
rect 27390 188852 46350 191312
rect 24930 188846 27388 188852
rect 43890 184967 46350 188852
rect 24633 182507 24639 184967
rect 27099 182507 46350 184967
rect -800 172888 1660 177688
rect -800 165348 1660 167688
rect 43890 165348 46350 182507
rect 582340 181430 584800 186230
rect -800 162888 3213 165348
rect 39658 162888 46350 165348
rect 151670 160310 162410 160340
rect 151670 158440 151710 160310
rect 162360 159780 162410 160310
rect 162360 159600 164610 159780
rect 162360 158440 162410 159600
rect 151670 158410 162410 158440
rect -800 124776 480 124888
rect 34270 124590 34710 124630
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect 34270 120160 34290 124590
rect -800 120048 480 120160
rect 34240 119850 34290 120160
rect 34180 119700 34290 119850
rect 34680 120160 34710 124590
rect 34680 119850 34770 120160
rect 34680 119700 34820 119850
rect 34180 119290 34820 119700
rect -800 118866 480 118978
rect 164430 118440 164610 159600
rect 184220 153700 184230 153705
rect 184220 153583 184225 153700
rect 184220 153578 184230 153583
rect 184347 153578 184353 153705
rect 192699 152355 192876 152361
rect 180376 152319 180541 152325
rect 192699 152183 192704 152188
rect 192871 152183 192876 152188
rect 192699 152178 192876 152183
rect 180376 152159 180381 152164
rect 180536 152159 180541 152164
rect 180376 152154 180541 152159
rect 582340 146830 584800 151630
rect 195081 146733 195193 146739
rect 185356 146689 185485 146695
rect 195081 146626 195086 146631
rect 195188 146626 195193 146631
rect 195081 146621 195193 146626
rect 185356 146565 185361 146570
rect 185480 146565 185485 146570
rect 185356 146560 185485 146565
rect 182348 145682 182492 145688
rect 182348 145543 182353 145548
rect 182487 145543 182492 145548
rect 182348 145538 182492 145543
rect 197430 141875 197770 141910
rect 185936 141841 186064 141847
rect 185936 141718 185941 141723
rect 186059 141718 186064 141723
rect 185936 141713 186064 141718
rect 197430 141805 197545 141875
rect 197609 141870 197770 141875
rect 197610 141810 197770 141870
rect 197609 141805 197770 141810
rect 197430 141700 197770 141805
rect 182679 141215 182852 141221
rect 182679 141047 182684 141052
rect 182847 141047 182852 141052
rect 182679 141042 182852 141047
rect 200910 136765 201330 136930
rect 582340 136830 584800 141630
rect 200910 136701 201065 136765
rect 201135 136701 201330 136765
rect 200910 136700 201070 136701
rect 201130 136700 201330 136701
rect 186760 136378 186938 136415
rect 186760 136314 186806 136378
rect 186876 136314 186938 136378
rect 186760 136313 186811 136314
rect 186871 136313 186938 136314
rect 186760 136267 186938 136313
rect 182943 135997 183150 136003
rect 200910 135940 201330 136700
rect 182943 135795 182948 135800
rect 183145 135795 183150 135800
rect 182943 135790 183150 135795
rect 171150 130045 171330 130070
rect 171150 129975 171195 130045
rect 171259 130040 171330 130045
rect 171260 129980 171330 130040
rect 171259 129975 171330 129980
rect 171150 129920 171330 129975
rect 205210 128370 205330 128390
rect 187089 128332 187201 128338
rect 205210 128310 205240 128370
rect 205300 128310 205330 128370
rect 205210 128270 205330 128310
rect 187089 128225 187094 128230
rect 187196 128225 187201 128230
rect 187089 128220 187201 128225
rect 183117 127744 183284 127750
rect 183117 127582 183122 127587
rect 183279 127582 183284 127587
rect 183117 127577 183284 127582
rect 206240 124455 206420 124500
rect 206240 124391 206305 124455
rect 206375 124391 206420 124455
rect 206240 124390 206310 124391
rect 206370 124390 206420 124391
rect 206240 124320 206420 124390
rect 183348 123805 183466 123811
rect 183348 123692 183353 123697
rect 183461 123692 183466 123697
rect 183348 123687 183466 123692
rect 187299 123741 187435 123756
rect 187299 123658 187321 123741
rect 187414 123658 187435 123741
rect 187299 123653 187326 123658
rect 187409 123653 187435 123658
rect 187299 123624 187435 123653
rect 187562 120886 187678 120892
rect 187562 120775 187567 120780
rect 187673 120775 187678 120780
rect 187562 120770 187678 120775
rect 207990 120765 208140 120810
rect 207990 120701 208015 120765
rect 208085 120701 208140 120765
rect 207990 120700 208020 120701
rect 208080 120700 208140 120701
rect 207990 120650 208140 120700
rect 183564 120064 183706 120070
rect 183564 119927 183569 119932
rect 183701 119927 183706 119932
rect 183564 119922 183706 119927
rect 164040 118260 181810 118440
rect 181030 113700 181430 113706
rect 180216 112195 180606 112201
rect 13584 103810 13590 103990
rect 13770 103810 14790 103990
rect 14610 102463 14790 103810
rect 180216 103749 180606 111805
rect 181030 103749 181430 113300
rect 180216 103351 180251 103749
rect 180649 103351 180655 103749
rect 181025 103351 181031 103749
rect 181429 103351 181435 103749
rect 180216 103094 180606 103351
rect 181030 103350 181430 103351
rect 180211 102706 180217 103094
rect 180605 102706 180611 103094
rect 180216 102705 180606 102706
rect 181630 102523 181810 118260
rect 184245 117491 184375 117497
rect 184245 117366 184250 117371
rect 184370 117366 184375 117371
rect 184245 117361 184375 117366
rect 187786 117396 188249 117533
rect 187786 117332 187971 117396
rect 188041 117332 188249 117396
rect 187786 117331 187976 117332
rect 188036 117331 188249 117332
rect 187786 117153 188249 117331
rect 187680 114460 188080 114466
rect 184250 114300 184650 114306
rect 182732 104274 182798 104279
rect 182732 104218 182737 104274
rect 182793 104218 182798 104274
rect 182732 104213 182798 104218
rect 182297 104038 182363 104043
rect 182297 103982 182302 104038
rect 182358 103982 182363 104038
rect 182297 103977 182363 103982
rect 182300 103204 182360 103977
rect 182735 103581 182795 104213
rect 183167 103962 183233 103967
rect 183167 103906 183172 103962
rect 183228 103906 183233 103962
rect 183167 103901 183233 103906
rect 182727 103517 182733 103581
rect 182797 103517 182803 103581
rect 183170 103213 183230 103901
rect 184250 103749 184650 113900
rect 185732 104890 185798 104895
rect 185732 104834 185737 104890
rect 185793 104834 185798 104890
rect 185732 104829 185798 104834
rect 185735 104612 185795 104829
rect 185727 104548 185733 104612
rect 185797 104548 185803 104612
rect 186168 104201 186232 104207
rect 186427 104199 186493 104202
rect 186232 104197 186493 104199
rect 186232 104141 186432 104197
rect 186488 104141 186493 104197
rect 186232 104139 186493 104141
rect 186168 104131 186232 104137
rect 186427 104136 186493 104139
rect 186586 103802 186684 103807
rect 186585 103801 186685 103802
rect 183602 103587 183668 103592
rect 183602 103531 183607 103587
rect 183663 103531 183668 103587
rect 182292 103140 182298 103204
rect 182362 103140 182368 103204
rect 183162 103149 183168 103213
rect 183232 103149 183238 103213
rect 183602 103172 183668 103531
rect 184245 103351 184251 103749
rect 184649 103351 184655 103749
rect 186585 103703 186586 103801
rect 186684 103703 186685 103801
rect 187680 103749 188080 114060
rect 190630 114230 191030 114236
rect 190630 106949 191030 113830
rect 190625 106551 190631 106949
rect 191029 106551 191035 106949
rect 190630 106550 191030 106551
rect 212340 105825 212940 106250
rect 212340 105761 212525 105825
rect 212595 105761 212940 105825
rect 212340 105760 212530 105761
rect 212590 105760 212940 105761
rect 212340 105440 212940 105760
rect 188733 104762 188797 104768
rect 192837 104760 192903 104763
rect 188797 104758 192903 104760
rect 188797 104702 192842 104758
rect 192898 104702 192903 104758
rect 188797 104700 192903 104702
rect 188733 104692 188797 104698
rect 192837 104697 192903 104700
rect 191483 104568 191549 104573
rect 191483 104512 191488 104568
rect 191544 104512 191549 104568
rect 191483 104507 191549 104512
rect 189090 104132 189290 104170
rect 189090 104068 189168 104132
rect 189232 104068 189290 104132
rect 189090 103980 189290 104068
rect 186585 103702 186685 103703
rect 186586 103697 186684 103702
rect 185297 103639 185363 103644
rect 185297 103583 185302 103639
rect 185358 103583 185363 103639
rect 185297 103578 185363 103583
rect 184250 103350 184650 103351
rect 185300 103178 185360 103578
rect 187675 103351 187681 103749
rect 188079 103351 188085 103749
rect 188281 103702 188381 103722
rect 188281 103638 188298 103702
rect 188362 103638 188381 103702
rect 188281 103620 188381 103638
rect 187680 103350 188080 103351
rect 183597 103108 183603 103172
rect 183667 103108 183673 103172
rect 185292 103114 185298 103178
rect 185362 103114 185368 103178
rect 189570 103142 189690 103170
rect 183602 103107 183668 103108
rect 189570 103078 189603 103142
rect 189667 103078 189690 103142
rect 189570 103030 189690 103078
rect 14560 102283 181070 102463
rect 191486 102382 191546 104507
rect 191478 102318 191484 102382
rect 191548 102318 191554 102382
rect 5790 102223 5970 102229
rect 5970 102043 181066 102223
rect 5790 102037 5970 102043
rect 192142 99387 192512 99392
rect 192141 99386 198982 99387
rect 192141 99016 192142 99386
rect 192512 99016 198982 99386
rect 192141 99015 198982 99016
rect 199354 99015 199360 99387
rect 192142 99010 192512 99015
rect 192142 98387 192512 98392
rect 192141 98386 198982 98387
rect 192141 98016 192142 98386
rect 192512 98016 198982 98386
rect 192141 98015 198982 98016
rect 199354 98015 199360 98387
rect 192142 98010 192512 98015
rect 192142 96387 192512 96392
rect 192141 96386 198982 96387
rect 192141 96016 192142 96386
rect 192512 96016 198982 96386
rect 192141 96015 198982 96016
rect 199354 96015 199360 96387
rect 192142 96010 192512 96015
rect 192142 95387 192512 95392
rect 192141 95386 198982 95387
rect 192141 95016 192142 95386
rect 192512 95016 198982 95386
rect 192141 95015 198982 95016
rect 199354 95015 199360 95387
rect 583520 95118 584800 95230
rect 192142 95010 192512 95015
rect 583520 93936 584800 94048
rect 192142 93387 192512 93392
rect 192141 93386 198982 93387
rect 192141 93016 192142 93386
rect 192512 93016 198982 93386
rect 192141 93015 198982 93016
rect 199354 93015 199360 93387
rect 192142 93010 192512 93015
rect 583520 92754 584800 92866
rect 10245 92695 10395 92701
rect 10245 92550 10250 92555
rect 10390 92550 10395 92555
rect 10245 92545 10395 92550
rect 192142 92387 192512 92392
rect 192141 92386 198982 92387
rect 192141 92016 192142 92386
rect 192512 92016 198982 92386
rect 192141 92015 198982 92016
rect 199354 92015 199360 92387
rect 192142 92010 192512 92015
rect 180439 91635 180445 91855
rect 180655 91850 180665 91855
rect 180660 91640 180665 91850
rect 180655 91635 180665 91640
rect 190900 91850 190910 91855
rect 190900 91640 190905 91850
rect 190900 91635 190910 91640
rect 191120 91635 191126 91855
rect 583520 91572 584800 91684
rect 143724 88783 143836 89496
rect 143724 88713 189775 88783
rect 143724 83976 143836 88713
rect 157172 88401 157178 88465
rect 157242 88463 157248 88465
rect 157242 88403 189800 88463
rect 157242 88401 157248 88403
rect 166143 87955 166149 88278
rect 166462 88273 166472 88278
rect 166467 87960 166472 88273
rect 202750 88270 202760 88275
rect 181887 87961 181893 88025
rect 181957 87961 181963 88025
rect 184887 87961 184893 88025
rect 184957 87961 184963 88025
rect 187887 87961 187893 88025
rect 187957 87961 187963 88025
rect 166462 87955 166472 87960
rect 181207 87698 181213 87762
rect 181277 87698 181283 87762
rect 22914 83864 143836 83976
rect -800 81661 4286 81666
rect -800 81559 4179 81661
rect 4281 81559 4286 81661
rect -800 81554 4286 81559
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect -800 38439 1886 38444
rect -800 38337 1779 38439
rect 1881 38337 1886 38439
rect -800 38332 1886 38337
rect 22914 37646 23026 83864
rect 179340 78170 179780 78290
rect 179340 78090 179500 78170
rect 179570 78165 179780 78170
rect 179575 78095 179780 78165
rect 179570 78090 179780 78095
rect 179340 77910 179780 78090
rect 7414 37534 23026 37646
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 7414 17022 7526 37534
rect 157725 29466 157847 29471
rect 157725 29450 157730 29466
rect 157570 29390 157730 29450
rect 157725 29354 157730 29390
rect 157842 29450 157847 29466
rect 181215 29450 181275 87698
rect 181547 87688 181553 87752
rect 181617 87688 181623 87752
rect 157842 29390 181275 29450
rect 157842 29354 157847 29390
rect 157725 29349 157847 29354
rect 181555 28720 181615 87688
rect 181895 79783 181955 87961
rect 182227 86998 182233 87062
rect 182297 86998 182303 87062
rect 182567 87008 182573 87072
rect 182637 87008 182643 87072
rect 181892 79778 181958 79783
rect 181892 79722 181897 79778
rect 181953 79722 181958 79778
rect 181892 79717 181958 79722
rect 182235 79693 182295 86998
rect 182232 79688 182298 79693
rect 182232 79632 182237 79688
rect 182293 79632 182298 79688
rect 182232 79627 182298 79632
rect 181930 78360 182320 78500
rect 181930 78355 182095 78360
rect 181930 78285 182090 78355
rect 181930 78280 182095 78285
rect 182165 78280 182320 78360
rect 181930 78110 182320 78280
rect 160750 28706 181615 28720
rect 160750 28660 161276 28706
rect 161271 28594 161276 28660
rect 161388 28660 181615 28706
rect 161388 28594 161393 28660
rect 161271 28589 161393 28594
rect 182575 27083 182635 87008
rect 182907 86978 182913 87042
rect 182977 86978 182983 87042
rect 183247 87008 183253 87072
rect 183317 87008 183323 87072
rect 183587 87038 183593 87102
rect 183657 87038 183663 87102
rect 182915 79983 182975 86978
rect 182912 79978 182978 79983
rect 182912 79922 182917 79978
rect 182973 79922 182978 79978
rect 182912 79917 182978 79922
rect 183255 79573 183315 87008
rect 183252 79568 183318 79573
rect 183252 79512 183257 79568
rect 183313 79512 183318 79568
rect 183252 79507 183318 79512
rect 182920 78245 183310 78380
rect 182920 78240 183090 78245
rect 183160 78240 183310 78245
rect 182920 78170 183085 78240
rect 183165 78170 183310 78240
rect 182920 77990 183310 78170
rect 182572 27078 182638 27083
rect 182572 27022 182577 27078
rect 182633 27022 182638 27078
rect 182572 27017 182638 27022
rect 182575 27000 182635 27017
rect 75680 26502 75850 26540
rect 75680 26438 75728 26502
rect 75792 26438 75850 26502
rect 75680 26390 75850 26438
rect 182547 23680 182669 23681
rect 183595 23680 183655 87038
rect 184215 80153 184275 87698
rect 184212 80148 184278 80153
rect 184212 80092 184217 80148
rect 184273 80092 184278 80148
rect 184212 80087 184278 80092
rect 184215 80060 184275 80087
rect 183870 78335 184370 78510
rect 183870 78330 184090 78335
rect 184160 78330 184370 78335
rect 183870 78260 184085 78330
rect 184165 78260 184370 78330
rect 183870 78060 184370 78260
rect 182480 23676 183655 23680
rect 182480 23620 182552 23676
rect 182547 23564 182552 23620
rect 182664 23620 183655 23676
rect 182664 23564 182669 23620
rect 182547 23559 182669 23564
rect -800 16910 7526 17022
rect -800 15728 480 15840
rect -800 14546 480 14658
rect -800 13364 480 13476
rect -800 12182 480 12294
rect -800 11000 480 11112
rect -800 9818 480 9930
rect -800 8636 480 8748
rect 69759 8651 69881 8657
rect 69759 8534 69764 8539
rect 69876 8534 69881 8539
rect 69759 8529 69881 8534
rect -800 7454 480 7566
rect 66359 7091 66481 7097
rect 66359 6974 66364 6979
rect 66476 6974 66481 6979
rect 66359 6969 66481 6974
rect -800 6272 480 6384
rect 62869 5711 62991 5717
rect 62869 5594 62874 5599
rect 62986 5594 62991 5599
rect 62869 5589 62991 5594
rect -800 5090 480 5202
rect 55239 4381 55361 4387
rect 55239 4264 55244 4269
rect 55356 4264 55361 4269
rect 55239 4259 55361 4264
rect -800 3908 480 4020
rect 52329 3351 52451 3357
rect 52329 3234 52334 3239
rect 52446 3234 52451 3239
rect 52329 3229 52451 3234
rect -800 2726 480 2838
rect 184555 2503 184615 87688
rect 184895 79783 184955 87961
rect 185227 86998 185233 87062
rect 185297 86998 185303 87062
rect 185567 87008 185573 87072
rect 185637 87008 185643 87072
rect 184892 79778 184958 79783
rect 184892 79722 184897 79778
rect 184953 79722 184958 79778
rect 184892 79717 184958 79722
rect 185235 79693 185295 86998
rect 185232 79688 185298 79693
rect 185232 79632 185237 79688
rect 185293 79632 185298 79688
rect 185232 79627 185298 79632
rect 184900 78165 185400 78340
rect 184900 78160 185090 78165
rect 185160 78160 185400 78165
rect 184900 78090 185085 78160
rect 185165 78090 185400 78160
rect 184900 77890 185400 78090
rect 185575 4453 185635 87008
rect 185907 86978 185913 87042
rect 185977 86978 185983 87042
rect 186247 87008 186253 87072
rect 186317 87008 186323 87072
rect 186587 87038 186593 87102
rect 186657 87038 186663 87102
rect 185915 79983 185975 86978
rect 185912 79978 185978 79983
rect 185912 79922 185917 79978
rect 185973 79922 185978 79978
rect 185912 79917 185978 79922
rect 186255 79573 186315 87008
rect 186252 79568 186318 79573
rect 186252 79512 186257 79568
rect 186313 79512 186318 79568
rect 186252 79507 186318 79512
rect 185920 78545 186330 78720
rect 185920 78540 186090 78545
rect 186160 78540 186330 78545
rect 185920 78470 186085 78540
rect 186165 78470 186330 78540
rect 185920 78300 186330 78470
rect 186595 6360 186655 87038
rect 187215 80153 187275 87698
rect 187212 80148 187278 80153
rect 187212 80092 187217 80148
rect 187273 80092 187278 80148
rect 187212 80087 187278 80092
rect 187215 80060 187275 80087
rect 186910 78655 187320 78840
rect 186910 78650 187090 78655
rect 187160 78650 187320 78655
rect 186910 78580 187085 78650
rect 187165 78580 187320 78650
rect 186910 78420 187320 78580
rect 187555 7280 187615 87688
rect 187895 79783 187955 87961
rect 202750 87960 202755 88270
rect 202750 87955 202760 87960
rect 203070 87955 203076 88275
rect 189587 87728 189593 87792
rect 189657 87728 189663 87792
rect 189595 87102 189655 87728
rect 188227 86998 188233 87062
rect 188297 86998 188303 87062
rect 188567 87008 188573 87072
rect 188637 87008 188643 87072
rect 187892 79778 187958 79783
rect 187892 79722 187897 79778
rect 187953 79722 187958 79778
rect 187892 79717 187958 79722
rect 188235 79693 188295 86998
rect 188232 79688 188298 79693
rect 188232 79632 188237 79688
rect 188293 79632 188298 79688
rect 188232 79627 188298 79632
rect 187920 78325 188330 78510
rect 187920 78320 188090 78325
rect 188160 78320 188330 78325
rect 187920 78250 188085 78320
rect 188165 78250 188330 78320
rect 187920 78090 188330 78250
rect 188575 8943 188635 87008
rect 188907 86978 188913 87042
rect 188977 86978 188983 87042
rect 189247 87008 189253 87072
rect 189317 87008 189323 87072
rect 189587 87038 189593 87102
rect 189657 87038 189663 87102
rect 188915 79983 188975 86978
rect 188912 79978 188978 79983
rect 188912 79922 188917 79978
rect 188973 79922 188978 79978
rect 188912 79917 188978 79922
rect 189255 79573 189315 87008
rect 189252 79568 189318 79573
rect 189252 79512 189257 79568
rect 189313 79512 189318 79568
rect 189252 79507 189318 79512
rect 188920 78495 189330 78650
rect 188920 78490 189090 78495
rect 189160 78490 189330 78495
rect 188920 78420 189085 78490
rect 189165 78420 189330 78490
rect 188920 78230 189330 78420
rect 189595 9750 189655 87038
rect 189930 78435 190340 78590
rect 189930 78430 190090 78435
rect 190160 78430 190340 78435
rect 189930 78360 190085 78430
rect 190165 78360 190340 78430
rect 189930 78170 190340 78360
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect 583520 16910 584800 17022
rect 583520 15728 584800 15840
rect 583520 14546 584800 14658
rect 583520 13364 584800 13476
rect 583520 12182 584800 12294
rect 583520 11000 584800 11112
rect 551331 10581 551453 10587
rect 551331 10464 551336 10469
rect 551448 10464 551453 10469
rect 551331 10459 551453 10464
rect 583520 9818 584800 9930
rect 239283 9806 239405 9811
rect 238164 9750 239288 9806
rect 189595 9694 239288 9750
rect 239400 9694 239405 9806
rect 189595 9690 239220 9694
rect 239283 9689 239405 9694
rect 576153 9741 576275 9747
rect 576153 9624 576158 9629
rect 576270 9624 576275 9629
rect 576153 9619 576275 9624
rect 188572 8938 188638 8943
rect 188572 8882 188577 8938
rect 188633 8882 188638 8938
rect 188572 8877 188638 8882
rect 583520 8636 584800 8748
rect 558423 7881 558545 7887
rect 558423 7764 558428 7769
rect 558540 7764 558545 7769
rect 558423 7759 558545 7764
rect 583520 7454 584800 7566
rect 218007 7286 218129 7291
rect 218007 7280 218012 7286
rect 187555 7220 218012 7280
rect 218007 7174 218012 7220
rect 218124 7280 218129 7286
rect 218124 7220 218530 7280
rect 218124 7174 218129 7220
rect 218007 7169 218129 7174
rect 572607 6561 572729 6567
rect 572607 6444 572612 6449
rect 572724 6444 572729 6449
rect 572607 6439 572729 6444
rect 210957 6360 211023 6363
rect 186595 6358 211023 6360
rect 186595 6302 210962 6358
rect 211018 6302 211023 6358
rect 186595 6300 211023 6302
rect 210957 6297 211023 6300
rect 565515 6311 565637 6317
rect 565515 6194 565520 6199
rect 565632 6194 565637 6199
rect 565515 6189 565637 6194
rect 569061 6291 569183 6297
rect 583520 6272 584800 6384
rect 569061 6174 569066 6179
rect 569178 6174 569183 6179
rect 569061 6169 569183 6174
rect 554877 6161 554999 6167
rect 554877 6044 554882 6049
rect 554994 6044 554999 6049
rect 554877 6039 554999 6044
rect 561969 6081 562091 6087
rect 561969 5964 561974 5969
rect 562086 5964 562091 5969
rect 561969 5959 562091 5964
rect 583520 5090 584800 5202
rect 185572 4448 185638 4453
rect 185572 4392 185577 4448
rect 185633 4392 185638 4448
rect 185572 4387 185638 4392
rect 583520 3908 584800 4020
rect 583520 2726 584800 2838
rect 184552 2498 184618 2503
rect 184552 2442 184557 2498
rect 184613 2442 184618 2498
rect 184552 2437 184618 2442
rect 49529 2271 49651 2277
rect 49529 2154 49534 2159
rect 49646 2154 49651 2159
rect 49529 2149 49651 2154
rect 46409 1731 46531 1737
rect -800 1544 480 1656
rect 46409 1614 46414 1619
rect 46526 1614 46531 1619
rect 46409 1609 46531 1614
rect 583520 1544 584800 1656
<< via3 >>
rect 22590 695320 23050 695780
rect 23590 695310 24050 695770
rect 24590 695420 25050 695880
rect 25590 695420 26050 695880
rect 165595 699685 168093 699689
rect 10251 683795 10389 683799
rect 10251 683665 10255 683795
rect 10255 683665 10385 683795
rect 10385 683665 10389 683795
rect 10251 683661 10389 683665
rect 165595 697195 165599 699685
rect 165599 697195 168089 699685
rect 168089 697195 168093 699685
rect 165595 697191 168093 697195
rect 218481 697631 220979 700129
rect 319171 698681 321669 701179
rect 26658 682328 26663 683627
rect 26663 682328 27687 683627
rect 27687 682328 27692 683627
rect 29711 682806 29716 683670
rect 29716 682806 30585 683670
rect 30585 682806 30590 683670
rect 31106 683151 31111 683644
rect 31111 683151 31609 683644
rect 31609 683151 31614 683644
rect 31106 683146 31614 683151
rect 29711 682801 30590 682806
rect 26658 682323 27692 682328
rect 22490 677810 24950 680270
rect 5721 673341 6039 673659
rect 14980 672355 15070 672360
rect 14980 672265 15065 672355
rect 15065 672265 15070 672355
rect 14980 672260 15070 672265
rect 19000 634750 21460 637210
rect 14060 559600 16520 562060
rect 14400 549750 16860 552210
rect 40191 689345 42649 689349
rect 40191 686895 40195 689345
rect 40195 686895 42645 689345
rect 42645 686895 42649 689345
rect 40191 686891 42649 686895
rect 569271 698981 569589 699299
rect 36783 295420 36895 295532
rect 29956 249971 30024 250039
rect 32588 206138 32652 206142
rect 32588 206082 32592 206138
rect 32592 206082 32648 206138
rect 32648 206082 32652 206138
rect 32588 206078 32652 206082
rect 24950 203217 26591 204858
rect 49575 204410 49645 204415
rect 49575 204351 49580 204410
rect 49580 204351 49640 204410
rect 49640 204351 49645 204410
rect 54111 211900 54175 211905
rect 54111 211840 54170 211900
rect 54170 211840 54175 211900
rect 54111 211835 54175 211840
rect 54510 209920 54574 209925
rect 54510 209860 54569 209920
rect 54569 209860 54574 209920
rect 54510 209855 54574 209860
rect 54945 207540 55009 207545
rect 54945 207480 55004 207540
rect 55004 207480 55009 207540
rect 54945 207475 55009 207480
rect 56525 205690 56595 205695
rect 56525 205631 56530 205690
rect 56530 205631 56590 205690
rect 56590 205631 56595 205690
rect 51752 202962 51816 203026
rect 53498 202998 53562 203002
rect 53498 202942 53502 202998
rect 53502 202942 53558 202998
rect 53558 202942 53562 202998
rect 53498 202938 53562 202942
rect 54838 202968 54902 202972
rect 54838 202912 54842 202968
rect 54842 202912 54898 202968
rect 54898 202912 54902 202968
rect 54838 202908 54902 202912
rect 55528 202948 55592 202952
rect 55528 202892 55532 202948
rect 55532 202892 55588 202948
rect 55588 202892 55592 202948
rect 55528 202888 55592 202892
rect 54227 202858 54291 202862
rect 54227 202802 54231 202858
rect 54231 202802 54287 202858
rect 54287 202802 54291 202858
rect 54227 202798 54291 202802
rect 44915 201070 45215 201075
rect 44915 200770 44920 201070
rect 44920 200770 45215 201070
rect 44915 200765 45215 200770
rect 24649 199640 25774 200765
rect 45015 200130 45315 200135
rect 45015 199830 45020 200130
rect 45020 199830 45315 200130
rect 45015 199825 45315 199830
rect 49184 199490 49254 199560
rect 45445 199110 45745 199115
rect 45445 198810 45450 199110
rect 45450 198810 45745 199110
rect 45445 198805 45745 198810
rect 24781 195324 27241 197784
rect 55765 196350 55865 196355
rect 55765 196250 55860 196350
rect 55860 196250 55865 196350
rect 55765 196245 55865 196250
rect 24930 188852 27390 191312
rect 24639 182507 27099 184967
rect 34290 119700 34680 124590
rect 184230 153700 184347 153705
rect 184230 153583 184342 153700
rect 184342 153583 184347 153700
rect 184230 153578 184347 153583
rect 192699 152350 192876 152355
rect 180376 152314 180541 152319
rect 180376 152164 180381 152314
rect 180381 152164 180536 152314
rect 180536 152164 180541 152314
rect 192699 152188 192704 152350
rect 192704 152188 192871 152350
rect 192871 152188 192876 152350
rect 195081 146728 195193 146733
rect 185356 146684 185485 146689
rect 185356 146570 185361 146684
rect 185361 146570 185480 146684
rect 185480 146570 185485 146684
rect 195081 146631 195086 146728
rect 195086 146631 195188 146728
rect 195188 146631 195193 146728
rect 182348 145677 182492 145682
rect 182348 145548 182353 145677
rect 182353 145548 182487 145677
rect 182487 145548 182492 145677
rect 185936 141836 186064 141841
rect 185936 141723 185941 141836
rect 185941 141723 186059 141836
rect 186059 141723 186064 141836
rect 197545 141870 197609 141875
rect 197545 141810 197550 141870
rect 197550 141810 197609 141870
rect 197545 141805 197609 141810
rect 182679 141210 182852 141215
rect 182679 141052 182684 141210
rect 182684 141052 182847 141210
rect 182847 141052 182852 141210
rect 201065 136760 201135 136765
rect 201065 136701 201070 136760
rect 201070 136701 201130 136760
rect 201130 136701 201135 136760
rect 186806 136373 186876 136378
rect 186806 136314 186811 136373
rect 186811 136314 186871 136373
rect 186871 136314 186876 136373
rect 182943 135992 183150 135997
rect 182943 135800 182948 135992
rect 182948 135800 183145 135992
rect 183145 135800 183150 135992
rect 171195 130040 171259 130045
rect 171195 129980 171200 130040
rect 171200 129980 171259 130040
rect 171195 129975 171259 129980
rect 187089 128327 187201 128332
rect 187089 128230 187094 128327
rect 187094 128230 187196 128327
rect 187196 128230 187201 128327
rect 183117 127739 183284 127744
rect 183117 127587 183122 127739
rect 183122 127587 183279 127739
rect 183279 127587 183284 127739
rect 206305 124450 206375 124455
rect 206305 124391 206310 124450
rect 206310 124391 206370 124450
rect 206370 124391 206375 124450
rect 183348 123800 183466 123805
rect 183348 123697 183353 123800
rect 183353 123697 183461 123800
rect 183461 123697 183466 123800
rect 187321 123736 187414 123741
rect 187321 123658 187326 123736
rect 187326 123658 187409 123736
rect 187409 123658 187414 123736
rect 187562 120881 187678 120886
rect 187562 120780 187567 120881
rect 187567 120780 187673 120881
rect 187673 120780 187678 120881
rect 208015 120760 208085 120765
rect 208015 120701 208020 120760
rect 208020 120701 208080 120760
rect 208080 120701 208085 120760
rect 183564 120059 183706 120064
rect 183564 119932 183569 120059
rect 183569 119932 183701 120059
rect 183701 119932 183706 120059
rect 181030 113300 181430 113700
rect 180216 111805 180606 112195
rect 13590 103810 13770 103990
rect 180251 103351 180649 103749
rect 181031 103351 181429 103749
rect 180217 102706 180605 103094
rect 184245 117486 184375 117491
rect 184245 117371 184250 117486
rect 184250 117371 184370 117486
rect 184370 117371 184375 117486
rect 187971 117391 188041 117396
rect 187971 117332 187976 117391
rect 187976 117332 188036 117391
rect 188036 117332 188041 117391
rect 184250 113900 184650 114300
rect 182733 103517 182797 103581
rect 187680 114060 188080 114460
rect 185733 104548 185797 104612
rect 186168 104137 186232 104201
rect 182298 103140 182362 103204
rect 183168 103149 183232 103213
rect 184251 103351 184649 103749
rect 186586 103797 186684 103801
rect 186586 103707 186590 103797
rect 186590 103707 186680 103797
rect 186680 103707 186684 103797
rect 186586 103703 186684 103707
rect 190630 113830 191030 114230
rect 190631 106551 191029 106949
rect 212525 105820 212595 105825
rect 212525 105761 212530 105820
rect 212530 105761 212590 105820
rect 212590 105761 212595 105820
rect 188733 104698 188797 104762
rect 189168 104128 189232 104132
rect 189168 104072 189172 104128
rect 189172 104072 189228 104128
rect 189228 104072 189232 104128
rect 189168 104068 189232 104072
rect 187681 103351 188079 103749
rect 188298 103698 188362 103702
rect 188298 103642 188302 103698
rect 188302 103642 188358 103698
rect 188358 103642 188362 103698
rect 188298 103638 188362 103642
rect 183603 103108 183667 103172
rect 185298 103114 185362 103178
rect 189603 103138 189667 103142
rect 189603 103082 189607 103138
rect 189607 103082 189663 103138
rect 189663 103082 189667 103138
rect 189603 103078 189667 103082
rect 191484 102318 191548 102382
rect 5790 102043 5970 102223
rect 192142 99016 192512 99386
rect 198982 99015 199354 99387
rect 192142 98016 192512 98386
rect 198982 98015 199354 98387
rect 192142 96016 192512 96386
rect 198982 96015 199354 96387
rect 192142 95016 192512 95386
rect 198982 95015 199354 95387
rect 192142 93016 192512 93386
rect 198982 93015 199354 93387
rect 10245 92690 10395 92695
rect 10245 92555 10250 92690
rect 10250 92555 10390 92690
rect 10390 92555 10395 92690
rect 192142 92016 192512 92386
rect 198982 92015 199354 92387
rect 180445 91850 180655 91855
rect 180445 91640 180450 91850
rect 180450 91640 180655 91850
rect 180445 91635 180655 91640
rect 190910 91850 191120 91855
rect 190910 91640 191115 91850
rect 191115 91640 191120 91850
rect 190910 91635 191120 91640
rect 157178 88401 157242 88465
rect 166149 88273 166462 88278
rect 166149 87960 166154 88273
rect 166154 87960 166462 88273
rect 202760 88270 203070 88275
rect 181893 87961 181957 88025
rect 184893 87961 184957 88025
rect 187893 87961 187957 88025
rect 166149 87955 166462 87960
rect 181213 87698 181277 87762
rect 179500 78165 179570 78170
rect 179500 78095 179505 78165
rect 179505 78095 179570 78165
rect 179500 78090 179570 78095
rect 181553 87688 181617 87752
rect 182233 86998 182297 87062
rect 182573 87008 182637 87072
rect 182095 78355 182165 78360
rect 182095 78285 182160 78355
rect 182160 78285 182165 78355
rect 182095 78280 182165 78285
rect 182913 86978 182977 87042
rect 183253 87008 183317 87072
rect 183593 87038 183657 87102
rect 183085 78175 183090 78240
rect 183090 78175 183160 78240
rect 183160 78175 183165 78240
rect 183085 78170 183165 78175
rect 75728 26498 75792 26502
rect 75728 26442 75732 26498
rect 75732 26442 75788 26498
rect 75788 26442 75792 26498
rect 75728 26438 75792 26442
rect 184085 78265 184090 78330
rect 184090 78265 184160 78330
rect 184160 78265 184165 78330
rect 184085 78260 184165 78265
rect 69759 8646 69881 8651
rect 69759 8539 69764 8646
rect 69764 8539 69876 8646
rect 69876 8539 69881 8646
rect 66359 7086 66481 7091
rect 66359 6979 66364 7086
rect 66364 6979 66476 7086
rect 66476 6979 66481 7086
rect 62869 5706 62991 5711
rect 62869 5599 62874 5706
rect 62874 5599 62986 5706
rect 62986 5599 62991 5706
rect 55239 4376 55361 4381
rect 55239 4269 55244 4376
rect 55244 4269 55356 4376
rect 55356 4269 55361 4376
rect 52329 3346 52451 3351
rect 52329 3239 52334 3346
rect 52334 3239 52446 3346
rect 52446 3239 52451 3346
rect 185233 86998 185297 87062
rect 185573 87008 185637 87072
rect 185085 78095 185090 78160
rect 185090 78095 185160 78160
rect 185160 78095 185165 78160
rect 185085 78090 185165 78095
rect 185913 86978 185977 87042
rect 186253 87008 186317 87072
rect 186593 87038 186657 87102
rect 186085 78475 186090 78540
rect 186090 78475 186160 78540
rect 186160 78475 186165 78540
rect 186085 78470 186165 78475
rect 187085 78585 187090 78650
rect 187090 78585 187160 78650
rect 187160 78585 187165 78650
rect 187085 78580 187165 78585
rect 202760 87960 203065 88270
rect 203065 87960 203070 88270
rect 202760 87955 203070 87960
rect 189593 87728 189657 87792
rect 188233 86998 188297 87062
rect 188573 87008 188637 87072
rect 188085 78255 188090 78320
rect 188090 78255 188160 78320
rect 188160 78255 188165 78320
rect 188085 78250 188165 78255
rect 188913 86978 188977 87042
rect 189253 87008 189317 87072
rect 189593 87038 189657 87102
rect 189085 78425 189090 78490
rect 189090 78425 189160 78490
rect 189160 78425 189165 78490
rect 189085 78420 189165 78425
rect 190085 78365 190090 78430
rect 190090 78365 190160 78430
rect 190160 78365 190165 78430
rect 190085 78360 190165 78365
rect 551331 10576 551453 10581
rect 551331 10469 551336 10576
rect 551336 10469 551448 10576
rect 551448 10469 551453 10576
rect 576153 9736 576275 9741
rect 576153 9629 576158 9736
rect 576158 9629 576270 9736
rect 576270 9629 576275 9736
rect 558423 7876 558545 7881
rect 558423 7769 558428 7876
rect 558428 7769 558540 7876
rect 558540 7769 558545 7876
rect 572607 6556 572729 6561
rect 572607 6449 572612 6556
rect 572612 6449 572724 6556
rect 572724 6449 572729 6556
rect 565515 6306 565637 6311
rect 565515 6199 565520 6306
rect 565520 6199 565632 6306
rect 565632 6199 565637 6306
rect 569061 6286 569183 6291
rect 569061 6179 569066 6286
rect 569066 6179 569178 6286
rect 569178 6179 569183 6286
rect 554877 6156 554999 6161
rect 554877 6049 554882 6156
rect 554882 6049 554994 6156
rect 554994 6049 554999 6156
rect 561969 6076 562091 6081
rect 561969 5969 561974 6076
rect 561974 5969 562086 6076
rect 562086 5969 562091 6076
rect 49529 2266 49651 2271
rect 49529 2159 49534 2266
rect 49534 2159 49646 2266
rect 49646 2159 49651 2266
rect 46409 1726 46531 1731
rect 46409 1619 46414 1726
rect 46414 1619 46526 1726
rect 46526 1619 46531 1726
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 165594 699689 168094 702300
rect 165594 697191 165595 699689
rect 168093 697191 168094 699689
rect 218480 700129 220980 702300
rect 218480 697631 218481 700129
rect 220979 697631 220980 700129
rect 218480 697630 220980 697631
rect 319170 701179 321670 702300
rect 319170 698681 319171 701179
rect 321669 698681 321670 701179
rect 569270 699299 569590 699300
rect 569270 698981 569271 699299
rect 569589 698981 569590 699299
rect 569270 698980 569590 698981
rect 165594 697190 168094 697191
rect 319170 696530 321670 698681
rect 23049 695780 23051 695781
rect 23050 695320 23051 695780
rect 23049 695319 23051 695320
rect 20970 691430 42990 693890
rect 20970 684190 23430 691430
rect 40190 690040 42650 691430
rect 35930 689349 42910 690040
rect 35930 686891 40191 689349
rect 42649 686891 42910 689349
rect 35930 686320 42910 686891
rect 40190 684190 42650 686320
rect 10250 683799 10390 683950
rect 10250 683661 10251 683799
rect 10389 683661 10390 683799
rect 5720 673659 6040 673660
rect 5720 673341 5721 673659
rect 6039 673341 6040 673659
rect 5720 673340 6040 673341
rect 10250 92696 10390 683661
rect 20970 683670 42650 684190
rect 20970 683627 29711 683670
rect 20970 682323 26658 683627
rect 27692 682801 29711 683627
rect 30590 683644 42650 683670
rect 30590 683146 31106 683644
rect 31614 683146 42650 683644
rect 30590 682801 42650 683146
rect 27692 682323 42650 682801
rect 20970 681730 42650 682323
rect 22489 680270 22491 680271
rect 22489 677810 22490 680270
rect 22489 677809 22491 677810
rect 14979 672360 15071 672361
rect 14979 672260 14980 672360
rect 15070 672355 15071 672360
rect 15070 672265 17160 672355
rect 15070 672260 15071 672265
rect 14979 672259 15071 672260
rect 18999 637210 19001 637211
rect 18999 634750 19000 637210
rect 18999 634749 19001 634750
rect 14059 562060 16521 562061
rect 36140 562060 38600 681730
rect 40190 562060 42650 681730
rect 14059 559600 14060 562060
rect 16520 559600 44190 562060
rect 14059 559599 16521 559600
rect 14399 552210 16861 552211
rect 24506 552210 26966 559600
rect 36140 552210 38600 559600
rect 14399 549750 14400 552210
rect 16860 549750 38600 552210
rect 14399 549749 16861 549750
rect 24506 204858 26966 549750
rect 36829 295533 36889 297140
rect 36782 295532 36896 295533
rect 36782 295420 36783 295532
rect 36895 295420 36896 295532
rect 36782 295419 36896 295420
rect 24506 203217 24950 204858
rect 26591 203217 26966 204858
rect 24506 200765 26966 203217
rect 24506 199640 24649 200765
rect 25774 199640 26966 200765
rect 24506 197785 26966 199640
rect 29955 250039 30025 250040
rect 29955 249971 29956 250039
rect 30024 249971 30025 250039
rect 29955 199560 30025 249971
rect 36829 209382 36889 295419
rect 36829 209322 50973 209382
rect 32587 206142 32653 206143
rect 32587 206078 32588 206142
rect 32652 206140 32653 206142
rect 49580 206140 49640 206350
rect 32652 206080 49640 206140
rect 32652 206078 32653 206080
rect 32587 206077 32653 206078
rect 49580 204416 49640 206080
rect 49574 204415 49646 204416
rect 49574 204351 49575 204415
rect 49645 204351 49646 204415
rect 49574 204350 49646 204351
rect 50913 202301 50973 209322
rect 53510 207580 53570 213020
rect 54020 210237 54080 210740
rect 54020 210177 54298 210237
rect 54020 210077 54080 210177
rect 54238 208290 54298 210177
rect 54211 208230 54479 208290
rect 54238 208223 54298 208230
rect 53984 207580 54044 207688
rect 53510 207520 54044 207580
rect 53510 207488 53570 207520
rect 53984 204790 54044 207520
rect 54419 204750 54479 208230
rect 54640 207000 54700 208520
rect 54640 206940 54914 207000
rect 54854 204750 54914 206940
rect 55289 204750 55349 206470
rect 51751 203026 51817 203027
rect 51751 202962 51752 203026
rect 51816 202962 51817 203026
rect 51751 202961 51817 202962
rect 53497 203002 53563 203003
rect 51754 202301 51814 202961
rect 53497 202938 53498 203002
rect 53562 203000 53563 203002
rect 53794 203000 53854 203130
rect 53562 202940 53854 203000
rect 53562 202938 53563 202940
rect 53497 202937 53563 202938
rect 54229 202863 54289 203120
rect 54664 202970 54724 203110
rect 54837 202972 54903 202973
rect 54837 202970 54838 202972
rect 54664 202910 54838 202970
rect 54837 202908 54838 202910
rect 54902 202908 54903 202972
rect 54837 202907 54903 202908
rect 55099 202950 55159 203110
rect 55527 202952 55593 202953
rect 55527 202950 55528 202952
rect 55099 202890 55528 202950
rect 55527 202888 55528 202890
rect 55592 202950 55593 202952
rect 55592 202890 55600 202950
rect 55592 202888 55593 202890
rect 55527 202887 55593 202888
rect 54226 202862 54292 202863
rect 54226 202798 54227 202862
rect 54291 202798 54292 202862
rect 54226 202797 54292 202798
rect 50913 202241 51814 202301
rect 44914 201075 45216 201076
rect 44914 200765 44915 201075
rect 45215 200765 45216 201075
rect 44914 200764 45216 200765
rect 45014 200135 45316 200136
rect 45014 199825 45015 200135
rect 45315 199825 45316 200135
rect 45014 199824 45316 199825
rect 49183 199560 49255 199561
rect 29955 199490 49184 199560
rect 49254 199490 49255 199560
rect 49183 199489 49255 199490
rect 45444 199115 45746 199116
rect 45444 198805 45445 199115
rect 45745 198805 45746 199115
rect 45444 198804 45746 198805
rect 24506 197784 27242 197785
rect 24506 195324 24781 197784
rect 27241 195324 27242 197784
rect 24506 195323 27242 195324
rect 24506 191313 26966 195323
rect 24506 191312 27391 191313
rect 24506 188852 24930 191312
rect 27390 188852 27391 191312
rect 24506 188851 27391 188852
rect 24506 184968 26966 188851
rect 24506 184967 27100 184968
rect 24506 182507 24639 184967
rect 27099 182507 27100 184967
rect 24506 182506 27100 182507
rect 24506 181365 26966 182506
rect 34190 124590 34820 124690
rect 34190 119850 34290 124590
rect 34180 119700 34290 119850
rect 34680 119700 34820 124590
rect 34180 119440 34300 119700
rect 34620 119440 34820 119700
rect 34180 119290 34820 119440
rect 10244 92695 10396 92696
rect 10244 92555 10245 92695
rect 10395 92555 10396 92695
rect 10244 92554 10396 92555
rect 46414 13050 46526 13066
rect 53050 13050 53110 198800
rect 45470 12990 53110 13050
rect 46414 1732 46526 12990
rect 49534 11770 49646 11956
rect 53390 11770 53450 198800
rect 48760 11710 53450 11770
rect 49534 2272 49646 11710
rect 52334 6940 52446 7926
rect 53730 6940 53790 198800
rect 54070 11260 54130 198800
rect 54410 15140 54470 198800
rect 54750 19490 54810 198800
rect 55090 25220 55150 198800
rect 55430 26500 55490 198800
rect 55764 196355 55866 196356
rect 55764 196245 55765 196355
rect 55865 196245 55866 196355
rect 55764 196244 55866 196245
rect 180381 153780 180536 153827
rect 177860 153705 250110 153780
rect 177860 153578 184230 153705
rect 184347 153578 250110 153705
rect 177860 153460 250110 153578
rect 180381 152320 180536 153460
rect 192704 152356 192871 153460
rect 192698 152355 192877 152356
rect 180375 152319 180542 152320
rect 180375 152164 180376 152319
rect 180541 152164 180542 152319
rect 192698 152188 192699 152355
rect 192876 152188 192877 152355
rect 192698 152187 192877 152188
rect 180375 152163 180542 152164
rect 176500 146733 242990 146840
rect 176500 146689 195081 146733
rect 176500 146570 185356 146689
rect 185485 146631 195081 146689
rect 195193 146631 242990 146733
rect 185485 146570 242990 146631
rect 176500 146520 242990 146570
rect 182353 145683 182487 146520
rect 182347 145682 182493 145683
rect 182347 145548 182348 145682
rect 182492 145548 182493 145682
rect 182347 145547 182493 145548
rect 178584 141875 237680 141910
rect 178584 141841 197545 141875
rect 178584 141723 185936 141841
rect 186064 141805 197545 141841
rect 197609 141805 237680 141875
rect 186064 141723 237680 141805
rect 178584 141590 237680 141723
rect 182684 141216 182847 141590
rect 182678 141215 182853 141216
rect 182678 141052 182679 141215
rect 182852 141052 182853 141215
rect 182678 141051 182853 141052
rect 200910 136765 201330 136920
rect 200910 136701 201065 136765
rect 201135 136701 201330 136765
rect 200910 136530 201330 136701
rect 182075 136378 231710 136530
rect 182075 136314 186806 136378
rect 186876 136314 231710 136378
rect 182075 136210 231710 136314
rect 182948 135998 183145 136210
rect 182942 135997 183151 135998
rect 182942 135800 182943 135997
rect 183150 135800 183151 135997
rect 200910 135940 201330 136210
rect 182942 135799 183151 135800
rect 182100 128332 224620 128450
rect 182100 128230 187089 128332
rect 187201 128230 224620 128332
rect 182100 128130 224620 128230
rect 183122 127745 183279 128130
rect 183116 127744 183285 127745
rect 183116 127587 183117 127744
rect 183284 127587 183285 127744
rect 183116 127586 183285 127587
rect 179300 124455 219270 124530
rect 179300 124391 206305 124455
rect 206375 124391 219270 124455
rect 179300 124210 219270 124391
rect 183353 123806 183461 124210
rect 183347 123805 183467 123806
rect 183347 123697 183348 123805
rect 183466 123697 183467 123805
rect 187326 123742 187409 124210
rect 183347 123696 183467 123697
rect 187320 123741 187415 123742
rect 187320 123658 187321 123741
rect 187414 123658 187415 123741
rect 187320 123657 187415 123658
rect 187561 120886 187679 120887
rect 187561 120880 187562 120886
rect 176990 120780 187562 120880
rect 187678 120880 187679 120886
rect 187678 120780 214260 120880
rect 176990 120765 214260 120780
rect 176990 120701 208015 120765
rect 208085 120701 214260 120765
rect 176990 120560 214260 120701
rect 183569 120065 183701 120560
rect 183563 120064 183707 120065
rect 183563 119932 183564 120064
rect 183706 119932 183707 120064
rect 183563 119931 183707 119932
rect 187679 114460 187681 114461
rect 187679 114060 187680 114460
rect 187679 114059 187681 114060
rect 184249 113900 184250 113901
rect 184650 113900 184651 113901
rect 184249 113899 184651 113900
rect 181029 113300 181030 113301
rect 181430 113300 181431 113301
rect 181029 113299 181431 113300
rect 180215 111805 180216 111806
rect 180606 111805 180607 111806
rect 180215 111804 180607 111805
rect 185830 106896 186230 113640
rect 185830 106544 185854 106896
rect 186206 106544 186230 106896
rect 189600 106976 190000 113390
rect 213940 110940 214260 120560
rect 218950 114550 219270 124210
rect 224300 116630 224620 128130
rect 231390 119390 231710 136210
rect 237360 121630 237680 141590
rect 242670 124620 242990 146520
rect 249790 131040 250110 153460
rect 249790 131016 576374 131040
rect 249790 130744 576078 131016
rect 576350 130744 576374 131016
rect 249790 130720 576374 130744
rect 242670 124596 572828 124620
rect 242670 124324 572532 124596
rect 572804 124324 572828 124596
rect 242670 124300 572828 124324
rect 237360 121606 569282 121630
rect 237360 121334 568986 121606
rect 569258 121334 569282 121606
rect 237360 121310 569282 121334
rect 231390 119366 565736 119390
rect 231390 119094 565440 119366
rect 565712 119094 565736 119366
rect 231390 119070 565736 119094
rect 224300 116606 562190 116630
rect 224300 116334 561894 116606
rect 562166 116334 562190 116606
rect 224300 116310 562190 116334
rect 218950 114526 558644 114550
rect 218950 114254 558348 114526
rect 558620 114254 558644 114526
rect 218950 114230 558644 114254
rect 213940 110916 555098 110940
rect 213940 110644 554802 110916
rect 555074 110644 555098 110916
rect 213940 110620 555098 110644
rect 189600 106624 189624 106976
rect 189976 106624 190000 106976
rect 189600 106600 190000 106624
rect 190630 106949 191030 106950
rect 190630 106551 190631 106949
rect 191029 106551 191030 106949
rect 190630 106550 191030 106551
rect 185830 106520 186230 106544
rect 174508 105159 196707 106225
rect 174508 91850 175574 105159
rect 188732 104762 188798 104763
rect 188732 104698 188733 104762
rect 188797 104698 188798 104762
rect 188732 104697 188798 104698
rect 185732 104612 185798 104613
rect 185732 104548 185733 104612
rect 185797 104548 185798 104612
rect 185732 104547 185798 104548
rect 180250 103749 180650 103750
rect 180250 103351 180251 103749
rect 180649 103351 180650 103749
rect 180250 103350 180650 103351
rect 181030 103749 181430 103750
rect 181030 103351 181031 103749
rect 181429 103351 181430 103749
rect 184250 103749 184650 103750
rect 182732 103581 182798 103582
rect 182732 103517 182733 103581
rect 182797 103517 182798 103581
rect 182732 103516 182798 103517
rect 181030 103350 181430 103351
rect 182297 103204 182363 103243
rect 182297 103140 182298 103204
rect 182362 103140 182363 103204
rect 182297 103139 182363 103140
rect 180216 103094 180606 103095
rect 180216 102706 180217 103094
rect 180605 102706 180606 103094
rect 182300 102710 182360 103139
rect 180216 101663 180606 102706
rect 182735 102703 182795 103516
rect 184250 103351 184251 103749
rect 184649 103351 184650 103749
rect 184250 103350 184650 103351
rect 183167 103213 183233 103214
rect 183167 103149 183168 103213
rect 183232 103149 183233 103213
rect 185297 103178 185363 103179
rect 183167 103148 183233 103149
rect 183602 103172 183668 103173
rect 183170 102733 183230 103148
rect 183602 103108 183603 103172
rect 183667 103108 183668 103172
rect 185297 103114 185298 103178
rect 185362 103114 185363 103178
rect 185297 103113 185363 103114
rect 183602 102695 183668 103108
rect 185300 102706 185360 103113
rect 185735 102697 185795 104547
rect 186167 104201 186233 104202
rect 186167 104137 186168 104201
rect 186232 104137 186233 104201
rect 186167 104136 186233 104137
rect 186170 102701 186230 104136
rect 186585 103801 186685 103802
rect 186585 103703 186586 103801
rect 186684 103703 186685 103801
rect 186585 103702 186685 103703
rect 187680 103749 188080 103750
rect 186605 102713 186665 103702
rect 187680 103351 187681 103749
rect 188079 103351 188080 103749
rect 188297 103702 188363 103703
rect 188297 103638 188298 103702
rect 188362 103638 188363 103702
rect 188297 103637 188363 103638
rect 187680 103350 188080 103351
rect 188300 102713 188360 103637
rect 188735 102690 188795 104697
rect 189167 104132 189233 104133
rect 189167 104068 189168 104132
rect 189232 104068 189233 104132
rect 189167 104067 189233 104068
rect 189170 102700 189230 104067
rect 189602 103142 189668 103143
rect 189602 103078 189603 103142
rect 189667 103078 189668 103142
rect 189602 103077 189668 103078
rect 189605 102690 189665 103077
rect 191483 102382 191549 102383
rect 191483 102318 191484 102382
rect 191548 102318 191549 102382
rect 191483 102317 191549 102318
rect 191486 101840 191546 102317
rect 195641 101309 196707 105159
rect 195641 100977 195986 101309
rect 196318 100977 196707 101309
rect 195641 100309 196707 100977
rect 195641 99977 195986 100309
rect 196318 99977 196707 100309
rect 192141 99386 192513 99387
rect 192141 99016 192142 99386
rect 192512 99016 192513 99386
rect 192141 99015 192513 99016
rect 195641 99309 196707 99977
rect 195641 98977 195986 99309
rect 196318 98977 196707 99309
rect 198981 99387 198983 99388
rect 198981 99015 198982 99387
rect 198981 99014 198983 99015
rect 192141 98386 192513 98387
rect 192141 98016 192142 98386
rect 192512 98016 192513 98386
rect 192141 98015 192513 98016
rect 195641 98309 196707 98977
rect 195641 97977 195986 98309
rect 196318 97977 196707 98309
rect 198981 98387 198983 98388
rect 198981 98015 198982 98387
rect 198981 98014 198983 98015
rect 195641 97309 196707 97977
rect 195641 96977 195986 97309
rect 196318 96977 196707 97309
rect 192141 96386 192513 96387
rect 192141 96016 192142 96386
rect 192512 96016 192513 96386
rect 192141 96015 192513 96016
rect 195641 96309 196707 96977
rect 195641 95977 195986 96309
rect 196318 95977 196707 96309
rect 198981 96387 198983 96388
rect 198981 96015 198982 96387
rect 198981 96014 198983 96015
rect 192141 95386 192513 95387
rect 192141 95016 192142 95386
rect 192512 95016 192513 95386
rect 192141 95015 192513 95016
rect 195641 95309 196707 95977
rect 195641 94977 195986 95309
rect 196318 94977 196707 95309
rect 198981 95387 198983 95388
rect 198981 95015 198982 95387
rect 198981 95014 198983 95015
rect 195641 94309 196707 94977
rect 195641 93977 195986 94309
rect 196318 93977 196707 94309
rect 192141 93386 192513 93387
rect 192141 93016 192142 93386
rect 192512 93016 192513 93386
rect 192141 93015 192513 93016
rect 195641 93309 196707 93977
rect 195641 92977 195986 93309
rect 196318 92977 196707 93309
rect 198981 93387 198983 93388
rect 198981 93015 198982 93387
rect 198981 93014 198983 93015
rect 192141 92386 192513 92387
rect 192141 92016 192142 92386
rect 192512 92016 192513 92386
rect 192141 92015 192513 92016
rect 195641 92309 196707 92977
rect 195641 91977 195986 92309
rect 196318 91977 196707 92309
rect 198981 92387 198983 92388
rect 198981 92015 198982 92387
rect 198981 92014 198983 92015
rect 180444 91855 180656 91856
rect 180444 91850 180445 91855
rect 174508 91640 180445 91850
rect 157177 88465 157243 88466
rect 157177 88463 157178 88465
rect 57480 88403 157178 88463
rect 157177 88401 157178 88403
rect 157242 88401 157243 88465
rect 157177 88400 157243 88401
rect 174508 86306 175574 91640
rect 176115 86306 176325 91640
rect 177115 86306 177325 91640
rect 178115 86306 178325 91640
rect 179115 86306 179325 91640
rect 180115 86306 180325 91640
rect 180444 91635 180445 91640
rect 180655 91635 180656 91855
rect 180444 91634 180656 91635
rect 190909 91855 191121 91856
rect 190909 91635 190910 91855
rect 191120 91850 191121 91855
rect 195641 91850 196707 91977
rect 191120 91640 196707 91850
rect 191120 91635 191145 91640
rect 190909 91634 191145 91635
rect 181892 88025 181958 88026
rect 181215 87763 181275 88023
rect 181212 87762 181278 87763
rect 181212 87698 181213 87762
rect 181277 87698 181278 87762
rect 181555 87753 181615 88023
rect 181892 87961 181893 88025
rect 181957 87961 181958 88025
rect 181892 87960 181958 87961
rect 181212 87697 181278 87698
rect 181552 87752 181618 87753
rect 181552 87688 181553 87752
rect 181617 87688 181618 87752
rect 181552 87687 181618 87688
rect 182235 87063 182295 88070
rect 182575 87073 182635 88080
rect 182572 87072 182638 87073
rect 182232 87062 182298 87063
rect 182232 86998 182233 87062
rect 182297 86998 182298 87062
rect 182572 87008 182573 87072
rect 182637 87008 182638 87072
rect 182915 87043 182975 88023
rect 183255 87073 183315 88023
rect 183595 87103 183655 88090
rect 184892 88025 184958 88026
rect 184892 87961 184893 88025
rect 184957 87961 184958 88025
rect 184892 87960 184958 87961
rect 183592 87102 183658 87103
rect 183252 87072 183318 87073
rect 182572 87007 182638 87008
rect 182912 87042 182978 87043
rect 182232 86997 182298 86998
rect 182912 86978 182913 87042
rect 182977 86978 182978 87042
rect 183252 87008 183253 87072
rect 183317 87008 183318 87072
rect 183592 87038 183593 87102
rect 183657 87038 183658 87102
rect 185235 87063 185295 88070
rect 185575 87073 185635 88080
rect 185572 87072 185638 87073
rect 183592 87037 183658 87038
rect 185232 87062 185298 87063
rect 183252 87007 183318 87008
rect 185232 86998 185233 87062
rect 185297 86998 185298 87062
rect 185572 87008 185573 87072
rect 185637 87008 185638 87072
rect 185915 87043 185975 88023
rect 186255 87073 186315 88023
rect 186595 87103 186655 88090
rect 187892 88025 187958 88026
rect 187892 87961 187893 88025
rect 187957 87961 187958 88025
rect 187892 87960 187958 87961
rect 186592 87102 186658 87103
rect 186252 87072 186318 87073
rect 185572 87007 185638 87008
rect 185912 87042 185978 87043
rect 185232 86997 185298 86998
rect 182912 86977 182978 86978
rect 185912 86978 185913 87042
rect 185977 86978 185978 87042
rect 186252 87008 186253 87072
rect 186317 87008 186318 87072
rect 186592 87038 186593 87102
rect 186657 87038 186658 87102
rect 188235 87063 188295 88070
rect 188575 87073 188635 88080
rect 188572 87072 188638 87073
rect 186592 87037 186658 87038
rect 188232 87062 188298 87063
rect 186252 87007 186318 87008
rect 188232 86998 188233 87062
rect 188297 86998 188298 87062
rect 188572 87008 188573 87072
rect 188637 87008 188638 87072
rect 188915 87043 188975 88023
rect 189255 87073 189315 88023
rect 189595 87793 189655 88100
rect 189592 87792 189658 87793
rect 189592 87728 189593 87792
rect 189657 87728 189658 87792
rect 189592 87727 189658 87728
rect 189595 87103 189655 87727
rect 189592 87102 189658 87103
rect 189252 87072 189318 87073
rect 188572 87007 188638 87008
rect 188912 87042 188978 87043
rect 188232 86997 188298 86998
rect 185912 86977 185978 86978
rect 188912 86978 188913 87042
rect 188977 86978 188978 87042
rect 189252 87008 189253 87072
rect 189317 87008 189318 87072
rect 189592 87038 189593 87102
rect 189657 87038 189658 87102
rect 189592 87037 189658 87038
rect 189252 87007 189318 87008
rect 188912 86977 188978 86978
rect 190935 86306 191145 91634
rect 191935 86306 192145 91640
rect 192935 86306 193145 91640
rect 193935 86306 194145 91640
rect 194935 86306 195145 91640
rect 195641 86306 196707 91640
rect 174119 85240 196707 86306
rect 174508 84804 175574 85240
rect 180287 84658 180610 84682
rect 180287 84383 180311 84658
rect 180586 84383 180610 84658
rect 180287 79182 180610 84383
rect 190631 84636 191030 84660
rect 190631 84285 190655 84636
rect 191006 84285 191030 84636
rect 190631 79010 191030 84285
rect 75727 26502 75793 26503
rect 75727 26500 75728 26502
rect 55430 26440 75728 26500
rect 75727 26438 75728 26440
rect 75792 26438 75793 26502
rect 75727 26437 75793 26438
rect 69764 25220 69876 25276
rect 55090 25160 70080 25220
rect 66364 19490 66476 19546
rect 54750 19430 67040 19490
rect 62874 15140 62986 15746
rect 54410 15080 63110 15140
rect 55244 11260 55356 11286
rect 54070 11200 58680 11260
rect 51770 6880 53790 6940
rect 52334 3352 52446 6880
rect 53730 6770 53790 6880
rect 55244 4382 55356 11200
rect 62874 5712 62986 15080
rect 66364 7092 66476 19430
rect 69764 8652 69876 25160
rect 69758 8651 69882 8652
rect 69758 8539 69759 8651
rect 69881 8539 69882 8651
rect 69758 8538 69882 8539
rect 66358 7091 66482 7092
rect 66358 6979 66359 7091
rect 66481 6979 66482 7091
rect 66358 6978 66482 6979
rect 62868 5711 62992 5712
rect 62868 5599 62869 5711
rect 62991 5599 62992 5711
rect 62868 5598 62992 5599
rect 55238 4381 55362 4382
rect 55238 4269 55239 4381
rect 55361 4269 55362 4381
rect 55238 4268 55362 4269
rect 52328 3351 52452 3352
rect 52328 3239 52329 3351
rect 52451 3239 52452 3351
rect 52328 3238 52452 3239
rect 49528 2271 49652 2272
rect 49528 2159 49529 2271
rect 49651 2159 49652 2271
rect 49528 2158 49652 2159
rect 46408 1731 46532 1732
rect 46408 1619 46409 1731
rect 46531 1619 46532 1731
rect 46408 1618 46532 1619
<< via4 >>
rect 569294 699004 569566 699276
rect 24589 695880 25051 695881
rect 22589 695780 23049 695781
rect 22589 695320 22590 695780
rect 22590 695320 23049 695780
rect 22589 695319 23049 695320
rect 23589 695770 24051 695771
rect 23589 695310 23590 695770
rect 23590 695310 24050 695770
rect 24050 695310 24051 695770
rect 24589 695420 24590 695880
rect 24590 695420 25050 695880
rect 25050 695420 25051 695880
rect 24589 695419 25051 695420
rect 25589 695880 26051 695881
rect 25589 695420 25590 695880
rect 25590 695420 26050 695880
rect 26050 695420 26051 695880
rect 25589 695419 26051 695420
rect 23589 695309 24051 695310
rect 5744 673364 6016 673636
rect 5720 102223 6040 102293
rect 5720 102043 5790 102223
rect 5790 102043 5970 102223
rect 5970 102043 6040 102223
rect 5720 101973 6040 102043
rect 22491 680270 24951 680271
rect 22491 677810 24950 680270
rect 24950 677810 24951 680270
rect 22491 677809 24951 677810
rect 17160 672150 17480 672470
rect 19001 637210 21461 637211
rect 19001 634750 21460 637210
rect 21460 634750 21461 637210
rect 19001 634749 21461 634750
rect 53380 213020 53700 213340
rect 53983 211905 54303 212030
rect 53983 211835 54111 211905
rect 54111 211835 54175 211905
rect 54175 211835 54303 211905
rect 53983 211710 54303 211835
rect 53890 210740 54210 211060
rect 54382 209925 54702 210050
rect 54382 209855 54510 209925
rect 54510 209855 54574 209925
rect 54574 209855 54702 209925
rect 54382 209730 54702 209855
rect 54510 208520 54830 208840
rect 54817 207545 55137 207670
rect 54817 207475 54945 207545
rect 54945 207475 55009 207545
rect 55009 207475 55137 207545
rect 54817 207350 55137 207475
rect 55159 206470 55479 206790
rect 56400 205695 56720 205823
rect 56400 205631 56525 205695
rect 56525 205631 56595 205695
rect 56595 205631 56720 205695
rect 56400 205503 56720 205631
rect 34300 119700 34620 119760
rect 34300 119440 34620 119700
rect 13520 103990 13840 104060
rect 13520 103810 13590 103990
rect 13590 103810 13770 103990
rect 13770 103810 13840 103990
rect 13520 103740 13840 103810
rect 171067 130045 171387 130170
rect 171067 129975 171195 130045
rect 171195 129975 171259 130045
rect 171259 129975 171387 130045
rect 171067 129850 171387 129975
rect 184150 117491 184470 117591
rect 184150 117371 184245 117491
rect 184245 117371 184375 117491
rect 184375 117371 184470 117491
rect 184150 117271 184470 117371
rect 187846 117396 188166 117524
rect 187846 117332 187971 117396
rect 187971 117332 188041 117396
rect 188041 117332 188166 117396
rect 187846 117204 188166 117332
rect 187681 114460 188081 114461
rect 184249 114300 184651 114301
rect 184249 113901 184250 114300
rect 184250 113901 184650 114300
rect 184650 113901 184651 114300
rect 187681 114060 188080 114460
rect 188080 114060 188081 114460
rect 187681 114059 188081 114060
rect 190629 114230 191031 114231
rect 181029 113700 181431 113701
rect 181029 113301 181030 113700
rect 181030 113301 181430 113700
rect 181430 113301 181431 113700
rect 185830 113640 186230 114040
rect 190629 113830 190630 114230
rect 190630 113830 191030 114230
rect 191030 113830 191031 114230
rect 190629 113829 191031 113830
rect 180215 112195 180607 112196
rect 180215 111806 180216 112195
rect 180216 111806 180606 112195
rect 180606 111806 180607 112195
rect 185854 106544 186206 106896
rect 189600 113390 190000 113790
rect 576078 130744 576350 131016
rect 572532 124324 572804 124596
rect 568986 121334 569258 121606
rect 565440 119094 565712 119366
rect 561894 116334 562166 116606
rect 558348 114254 558620 114526
rect 554802 110644 555074 110916
rect 189624 106624 189976 106976
rect 190654 106574 191006 106926
rect 212400 105825 212720 105953
rect 212400 105761 212525 105825
rect 212525 105761 212595 105825
rect 212595 105761 212720 105825
rect 212400 105633 212720 105761
rect 180274 103374 180626 103726
rect 181054 103374 181406 103726
rect 184274 103374 184626 103726
rect 187704 103374 188056 103726
rect 195986 100977 196318 101309
rect 195986 99977 196318 100309
rect 192165 99039 192489 99363
rect 195986 98977 196318 99309
rect 198983 99387 199355 99388
rect 198983 99015 199354 99387
rect 199354 99015 199355 99387
rect 198983 99014 199355 99015
rect 192165 98039 192489 98363
rect 195986 97977 196318 98309
rect 198983 98387 199355 98388
rect 198983 98015 199354 98387
rect 199354 98015 199355 98387
rect 198983 98014 199355 98015
rect 195986 96977 196318 97309
rect 192165 96039 192489 96363
rect 195986 95977 196318 96309
rect 198983 96387 199355 96388
rect 198983 96015 199354 96387
rect 199354 96015 199355 96387
rect 198983 96014 199355 96015
rect 192165 95039 192489 95363
rect 195986 94977 196318 95309
rect 198983 95387 199355 95388
rect 198983 95015 199354 95387
rect 199354 95015 199355 95387
rect 198983 95014 199355 95015
rect 195986 93977 196318 94309
rect 192165 93039 192489 93363
rect 195986 92977 196318 93309
rect 198983 93387 199355 93388
rect 198983 93015 199354 93387
rect 199354 93015 199355 93387
rect 198983 93014 199355 93015
rect 192165 92039 192489 92363
rect 195986 91977 196318 92309
rect 198983 92387 199355 92388
rect 198983 92015 199354 92387
rect 199354 92015 199355 92387
rect 198983 92014 199355 92015
rect 57160 88273 57480 88593
rect 166146 88278 166466 88279
rect 166146 87955 166149 88278
rect 166149 87955 166462 88278
rect 166462 87955 166466 88278
rect 166146 87954 166466 87955
rect 202755 88275 203075 88276
rect 202755 87955 202760 88275
rect 202760 87955 203070 88275
rect 203070 87955 203075 88275
rect 202755 87954 203075 87955
rect 180311 84383 180586 84658
rect 180287 78859 180610 79182
rect 190655 84285 191006 84636
rect 185965 78540 186285 78665
rect 181970 78360 182290 78480
rect 185965 78470 186085 78540
rect 186085 78470 186165 78540
rect 186165 78470 186285 78540
rect 179375 78170 179695 78290
rect 179375 78090 179500 78170
rect 179500 78090 179570 78170
rect 179570 78090 179695 78170
rect 181970 78280 182095 78360
rect 182095 78280 182165 78360
rect 182165 78280 182290 78360
rect 181970 78160 182290 78280
rect 182965 78240 183285 78365
rect 182965 78170 183085 78240
rect 183085 78170 183165 78240
rect 183165 78170 183285 78240
rect 179375 77970 179695 78090
rect 182965 78045 183285 78170
rect 183965 78330 184285 78455
rect 185965 78345 186285 78470
rect 186965 78650 187285 78775
rect 186965 78580 187085 78650
rect 187085 78580 187165 78650
rect 187165 78580 187285 78650
rect 186965 78455 187285 78580
rect 188965 78490 189285 78615
rect 190631 78611 191030 79010
rect 183965 78260 184085 78330
rect 184085 78260 184165 78330
rect 184165 78260 184285 78330
rect 187965 78320 188285 78445
rect 183965 78135 184285 78260
rect 184965 78160 185285 78285
rect 184965 78090 185085 78160
rect 185085 78090 185165 78160
rect 185165 78090 185285 78160
rect 187965 78250 188085 78320
rect 188085 78250 188165 78320
rect 188165 78250 188285 78320
rect 188965 78420 189085 78490
rect 189085 78420 189165 78490
rect 189165 78420 189285 78490
rect 188965 78295 189285 78420
rect 189965 78430 190285 78555
rect 189965 78360 190085 78430
rect 190085 78360 190165 78430
rect 190165 78360 190285 78430
rect 187965 78125 188285 78250
rect 189965 78235 190285 78360
rect 184965 77965 185285 78090
rect 551232 10581 551552 10685
rect 551232 10469 551331 10581
rect 551331 10469 551453 10581
rect 551453 10469 551552 10581
rect 551232 10365 551552 10469
rect 576054 9741 576374 9845
rect 576054 9629 576153 9741
rect 576153 9629 576275 9741
rect 576275 9629 576374 9741
rect 576054 9525 576374 9629
rect 558324 7881 558644 7985
rect 558324 7769 558423 7881
rect 558423 7769 558545 7881
rect 558545 7769 558644 7881
rect 558324 7665 558644 7769
rect 572508 6561 572828 6665
rect 572508 6449 572607 6561
rect 572607 6449 572729 6561
rect 572729 6449 572828 6561
rect 565416 6311 565736 6415
rect 554778 6161 555098 6265
rect 565416 6199 565515 6311
rect 565515 6199 565637 6311
rect 565637 6199 565736 6311
rect 554778 6049 554877 6161
rect 554877 6049 554999 6161
rect 554999 6049 555098 6161
rect 554778 5945 555098 6049
rect 561870 6081 562190 6185
rect 565416 6095 565736 6199
rect 568962 6291 569282 6395
rect 572508 6345 572828 6449
rect 568962 6179 569061 6291
rect 569061 6179 569183 6291
rect 569183 6179 569282 6291
rect 561870 5969 561969 6081
rect 561969 5969 562091 6081
rect 562091 5969 562190 6081
rect 568962 6075 569282 6179
rect 561870 5865 562190 5969
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 13570 699276 569670 699300
rect 13570 699004 569294 699276
rect 569566 699004 569670 699276
rect 13570 698980 569670 699004
rect 5720 673636 6040 674020
rect 5720 673364 5744 673636
rect 6016 673364 6040 673636
rect 5720 102317 6040 673364
rect 13570 104084 13890 698980
rect 16200 695881 52140 697010
rect 16200 695781 24589 695881
rect 16200 695319 22589 695781
rect 23049 695771 24589 695781
rect 23049 695319 23589 695771
rect 16200 695309 23589 695319
rect 24051 695419 24589 695771
rect 25051 695419 25589 695881
rect 26051 695419 52140 695881
rect 24051 695309 52140 695419
rect 16200 694550 52140 695309
rect 16200 680270 18660 694550
rect 22467 680271 24975 680295
rect 22467 680270 22491 680271
rect 16200 677830 22491 680270
rect 16300 677810 22491 677830
rect 22467 677809 22491 677810
rect 24951 680270 24975 680271
rect 49680 680270 52140 694550
rect 24951 677810 52140 680270
rect 24951 677809 25340 677810
rect 22467 677785 25340 677809
rect 17130 672494 17450 674430
rect 17130 672470 17504 672494
rect 17130 672150 17160 672470
rect 17480 672150 17504 672470
rect 17130 672126 17504 672150
rect 17130 130170 17450 672126
rect 18977 637211 21485 637235
rect 18977 634749 19001 637211
rect 21461 637210 21485 637211
rect 22880 637210 25340 677785
rect 26710 637210 29170 677810
rect 21461 634750 29170 637210
rect 21461 634749 21485 634750
rect 18977 634725 21485 634749
rect 336440 234570 336760 235580
rect 336400 234250 576374 234570
rect 53356 213340 53724 213364
rect 336440 213340 336760 234250
rect 53356 213020 53380 213340
rect 53700 213020 336760 213340
rect 338550 229440 338870 230130
rect 572508 229440 572828 231090
rect 338550 229120 572828 229440
rect 53356 212996 53724 213020
rect 53959 212030 54327 212054
rect 338550 212030 338870 229120
rect 53959 211710 53983 212030
rect 54303 211710 338870 212030
rect 340730 226010 341050 226430
rect 340730 225690 569282 226010
rect 53959 211686 54327 211710
rect 53866 211060 54234 211084
rect 340730 211060 341050 225690
rect 342450 223150 342770 223950
rect 342380 222830 565736 223150
rect 53866 210740 53890 211060
rect 54210 210740 341050 211060
rect 53866 210716 54234 210740
rect 54358 210050 54726 210074
rect 342450 210050 342770 222830
rect 344410 220290 344730 220460
rect 344380 219970 562190 220290
rect 54358 209730 54382 210050
rect 54702 209730 342770 210050
rect 54358 209706 54726 209730
rect 54486 208840 54854 208864
rect 344410 208840 344730 219970
rect 54486 208520 54510 208840
rect 54830 208520 344730 208840
rect 346240 215530 346560 215810
rect 346240 215210 558644 215530
rect 54486 208496 54854 208520
rect 54793 207670 55161 207694
rect 346240 207670 346560 215210
rect 554778 211080 555098 212500
rect 354950 210760 555098 211080
rect 54793 207350 54817 207670
rect 55137 207350 346560 207670
rect 54793 207326 55161 207350
rect 55135 206790 55503 206814
rect 355080 206790 355400 210760
rect 356420 208920 551552 209240
rect 55135 206470 55159 206790
rect 55479 206470 355400 206790
rect 55135 206446 55503 206470
rect 56400 206050 56720 206060
rect 356460 206050 356780 208920
rect 56400 206020 356780 206050
rect 56330 205823 356780 206020
rect 56330 205503 56400 205823
rect 56720 205730 356780 205823
rect 56720 205503 56940 205730
rect 56330 205460 56940 205503
rect 171043 130170 171411 130194
rect 17130 129850 171067 130170
rect 171387 129850 171411 130170
rect 171043 129826 171411 129850
rect 34276 119760 34644 119784
rect 34276 119440 34300 119760
rect 34620 119440 34644 119760
rect 34276 119416 34644 119440
rect 13496 104060 13890 104084
rect 13496 103740 13520 104060
rect 13840 103740 13890 104060
rect 13496 103716 13890 103740
rect 13570 103330 13890 103716
rect 5696 102293 6064 102317
rect 5696 101973 5720 102293
rect 6040 101973 6064 102293
rect 5696 101949 6064 101973
rect 34300 88593 34620 119416
rect 183296 117591 212150 117640
rect 183296 117320 184150 117591
rect 184126 117271 184150 117320
rect 184470 117524 212150 117591
rect 184470 117320 187846 117524
rect 184470 117271 184494 117320
rect 184126 117247 184494 117271
rect 187822 117204 187846 117320
rect 188166 117320 212150 117524
rect 188166 117204 188190 117320
rect 187822 117180 188190 117204
rect 165195 114461 204045 114995
rect 165195 114301 187681 114461
rect 165195 113901 184249 114301
rect 184651 114059 187681 114301
rect 188081 114231 204045 114461
rect 188081 114059 190629 114231
rect 184651 114040 190629 114059
rect 184651 113901 185830 114040
rect 165195 113701 185830 113901
rect 165195 113301 181029 113701
rect 181431 113640 185830 113701
rect 186230 113829 190629 114040
rect 191031 113829 204045 114231
rect 186230 113790 204045 113829
rect 186230 113640 189600 113790
rect 181431 113390 189600 113640
rect 190000 113390 204045 113790
rect 181431 113301 204045 113390
rect 165195 113165 204045 113301
rect 57136 88593 57504 88617
rect 32990 88273 57160 88593
rect 57480 88273 57504 88593
rect 34300 88180 34620 88273
rect 57136 88249 57504 88273
rect 165195 88279 167025 113165
rect 180216 112220 180606 113165
rect 180191 112196 180631 112220
rect 180191 111806 180215 112196
rect 180607 111806 180631 112196
rect 180191 111782 180631 111806
rect 165195 87954 166146 88279
rect 166466 87954 167025 88279
rect 165195 79360 167025 87954
rect 170665 107905 200365 109735
rect 170665 106408 172495 107905
rect 178850 106408 179170 107905
rect 191631 107185 192031 107905
rect 198535 107185 200365 107905
rect 189600 106976 190000 107000
rect 170665 106036 179170 106408
rect 170665 105408 172495 106036
rect 178850 105408 179170 106036
rect 170665 105036 179170 105408
rect 170665 104408 172495 105036
rect 178850 104408 179170 105036
rect 170665 104036 179170 104408
rect 170665 103408 172495 104036
rect 178850 103408 179170 104036
rect 185830 106896 186230 106920
rect 185830 106544 185854 106896
rect 186206 106544 186230 106896
rect 185830 103750 186230 106544
rect 189600 106624 189624 106976
rect 189976 106624 190000 106976
rect 189600 103750 190000 106624
rect 190630 106926 191030 106950
rect 190630 106574 190654 106926
rect 191006 106574 191030 106926
rect 190630 103750 191030 106574
rect 170665 103036 179170 103408
rect 180250 103726 191030 103750
rect 180250 103374 180274 103726
rect 180626 103374 181054 103726
rect 181406 103374 184274 103726
rect 184626 103374 187704 103726
rect 188056 103374 191030 103726
rect 180250 103350 191030 103374
rect 170665 102408 172495 103036
rect 178850 102408 179170 103036
rect 170665 102036 179170 102408
rect 170665 101408 172495 102036
rect 178850 101408 179170 102036
rect 170665 101036 179170 101408
rect 170665 100408 172495 101036
rect 178850 100408 179170 101036
rect 170665 100036 179170 100408
rect 170665 99408 172495 100036
rect 178850 99408 179170 100036
rect 170665 99036 179170 99408
rect 170665 98408 172495 99036
rect 178850 98408 179170 99036
rect 170665 98036 179170 98408
rect 170665 97408 172495 98036
rect 178850 97408 179170 98036
rect 170665 97036 179170 97408
rect 170665 96408 172495 97036
rect 178850 96408 179170 97036
rect 170665 96036 179170 96408
rect 170665 95408 172495 96036
rect 178850 95408 179170 96036
rect 170665 95036 179170 95408
rect 170665 94408 172495 95036
rect 178850 94408 179170 95036
rect 170665 94036 179170 94408
rect 170665 93408 172495 94036
rect 178850 93408 179170 94036
rect 170665 93036 179170 93408
rect 170665 92408 172495 93036
rect 178850 92408 179170 93036
rect 170665 92036 179170 92408
rect 180287 92270 180610 92433
rect 180220 92110 180610 92270
rect 170665 91408 172495 92036
rect 178850 91408 179170 92036
rect 170665 91036 179170 91408
rect 170665 90408 172495 91036
rect 178850 90408 179170 91036
rect 170665 90036 179170 90408
rect 170665 89408 172495 90036
rect 178850 89408 179170 90036
rect 170665 89036 179170 89408
rect 170665 88408 172495 89036
rect 178850 88408 179170 89036
rect 170665 88036 179170 88408
rect 170665 87408 172495 88036
rect 178850 87408 179170 88036
rect 170665 87036 179170 87408
rect 170665 86408 172495 87036
rect 178850 86408 179170 87036
rect 170665 86036 179170 86408
rect 170665 85408 172495 86036
rect 178850 85408 179170 86036
rect 170665 85036 179170 85408
rect 170665 83810 172495 85036
rect 178850 83810 179170 85036
rect 180287 84658 180610 92110
rect 190630 92000 191030 103350
rect 180287 84383 180311 84658
rect 180586 84383 180610 84658
rect 180287 84359 180610 84383
rect 190631 84636 191030 92000
rect 190631 84285 190655 84636
rect 191006 84285 191030 84636
rect 190631 84261 191030 84285
rect 191631 106785 200365 107185
rect 191631 104727 192031 106785
rect 198535 104727 200365 106785
rect 191631 104327 200365 104727
rect 191631 103411 192031 104327
rect 198535 103411 200365 104327
rect 191631 103011 200365 103411
rect 191631 99387 192031 103011
rect 195883 101333 196418 101445
rect 193286 101309 196418 101333
rect 193286 100977 195986 101309
rect 196318 100977 196418 101309
rect 193286 100953 196418 100977
rect 195883 100333 196418 100953
rect 193286 100309 196418 100333
rect 193286 99977 195986 100309
rect 196318 99977 196418 100309
rect 193286 99953 196418 99977
rect 191631 99363 192513 99387
rect 191631 99039 192165 99363
rect 192489 99039 192513 99363
rect 195883 99333 196418 99953
rect 191631 99015 192513 99039
rect 193286 99309 196418 99333
rect 191631 98387 192031 99015
rect 193286 98977 195986 99309
rect 196318 98977 196418 99309
rect 193286 98953 196418 98977
rect 191631 98363 192513 98387
rect 191631 98039 192165 98363
rect 192489 98039 192513 98363
rect 195883 98333 196418 98953
rect 191631 98015 192513 98039
rect 193286 98309 196418 98333
rect 191631 96387 192031 98015
rect 193286 97977 195986 98309
rect 196318 97977 196418 98309
rect 193286 97953 196418 97977
rect 195883 97333 196418 97953
rect 193286 97309 196418 97333
rect 193286 96977 195986 97309
rect 196318 96977 196418 97309
rect 193286 96953 196418 96977
rect 191631 96363 192513 96387
rect 191631 96039 192165 96363
rect 192489 96039 192513 96363
rect 195883 96333 196418 96953
rect 191631 96015 192513 96039
rect 193286 96309 196418 96333
rect 191631 95387 192031 96015
rect 193286 95977 195986 96309
rect 196318 95977 196418 96309
rect 193286 95953 196418 95977
rect 191631 95363 192513 95387
rect 191631 95039 192165 95363
rect 192489 95039 192513 95363
rect 195883 95333 196418 95953
rect 191631 95015 192513 95039
rect 193286 95309 196418 95333
rect 191631 93387 192031 95015
rect 193286 94977 195986 95309
rect 196318 94977 196418 95309
rect 193286 94953 196418 94977
rect 195883 94333 196418 94953
rect 193286 94309 196418 94333
rect 193286 93977 195986 94309
rect 196318 93977 196418 94309
rect 193286 93953 196418 93977
rect 191631 93363 192513 93387
rect 191631 93039 192165 93363
rect 192489 93039 192513 93363
rect 195883 93333 196418 93953
rect 191631 93015 192513 93039
rect 193286 93309 196418 93333
rect 191631 92387 192031 93015
rect 193286 92977 195986 93309
rect 196318 92977 196418 93309
rect 193286 92953 196418 92977
rect 191631 92363 192513 92387
rect 191631 92039 192165 92363
rect 192489 92039 192513 92363
rect 195883 92333 196418 92953
rect 191631 92015 192513 92039
rect 193286 92309 196418 92333
rect 191631 90375 192031 92015
rect 193286 91977 195986 92309
rect 196318 91977 196418 92309
rect 193286 91953 196418 91977
rect 195883 91848 196418 91953
rect 198535 99388 200365 103011
rect 198535 99014 198983 99388
rect 199355 99014 200365 99388
rect 198535 98388 200365 99014
rect 198535 98014 198983 98388
rect 199355 98014 200365 98388
rect 198535 96388 200365 98014
rect 198535 96014 198983 96388
rect 199355 96014 200365 96388
rect 198535 95388 200365 96014
rect 198535 95014 198983 95388
rect 199355 95014 200365 95388
rect 198535 93388 200365 95014
rect 198535 93014 198983 93388
rect 199355 93014 200365 93388
rect 198535 92388 200365 93014
rect 198535 92014 198983 92388
rect 199355 92014 200365 92388
rect 198535 90375 200365 92014
rect 191631 90003 200365 90375
rect 191631 89375 192031 90003
rect 198535 89375 200365 90003
rect 191631 89003 200365 89375
rect 191631 88375 192031 89003
rect 198535 88375 200365 89003
rect 191631 88003 200365 88375
rect 191631 87375 192031 88003
rect 198535 87375 200365 88003
rect 191631 87003 200365 87375
rect 191631 86375 192031 87003
rect 198535 86375 200365 87003
rect 191631 86003 200365 86375
rect 191631 85375 192031 86003
rect 198535 85375 200365 86003
rect 191631 85003 200365 85375
rect 191631 83810 192031 85003
rect 198535 83810 200365 85003
rect 170665 81980 200365 83810
rect 202215 88276 204045 113165
rect 211830 106020 212150 117320
rect 551232 106020 551552 208920
rect 211830 105953 551552 106020
rect 211830 105700 212400 105953
rect 212376 105633 212400 105700
rect 212720 105700 551552 105953
rect 212720 105633 212744 105700
rect 212376 105609 212744 105633
rect 202215 87954 202755 88276
rect 203075 87954 204045 88276
rect 170665 81395 172495 81980
rect 202215 79360 204045 87954
rect 165195 79182 204045 79360
rect 165195 78859 180287 79182
rect 180610 79010 204045 79182
rect 180610 78859 190631 79010
rect 165195 78775 190631 78859
rect 165195 78665 186965 78775
rect 165195 78480 185965 78665
rect 165195 78290 181970 78480
rect 165195 77970 179375 78290
rect 179695 78160 181970 78290
rect 182290 78455 185965 78480
rect 182290 78365 183965 78455
rect 182290 78160 182965 78365
rect 179695 78045 182965 78160
rect 183285 78135 183965 78365
rect 184285 78345 185965 78455
rect 186285 78455 186965 78665
rect 187285 78615 190631 78775
rect 187285 78455 188965 78615
rect 186285 78445 188965 78455
rect 186285 78345 187965 78445
rect 184285 78285 187965 78345
rect 184285 78135 184965 78285
rect 183285 78045 184965 78135
rect 179695 77970 184965 78045
rect 165195 77965 184965 77970
rect 185285 78125 187965 78285
rect 188285 78295 188965 78445
rect 189285 78611 190631 78615
rect 191030 78611 204045 79010
rect 189285 78555 204045 78611
rect 189285 78295 189965 78555
rect 188285 78235 189965 78295
rect 190285 78235 204045 78555
rect 188285 78125 204045 78235
rect 185285 77965 204045 78125
rect 165195 77530 204045 77965
rect 165195 75565 167025 77530
rect 551232 10709 551552 105700
rect 554778 110916 555098 210760
rect 554778 110644 554802 110916
rect 555074 110644 555098 110916
rect 551208 10685 551576 10709
rect 551208 10365 551232 10685
rect 551552 10365 551576 10685
rect 551208 10341 551576 10365
rect 554778 6289 555098 110644
rect 558324 114526 558644 215210
rect 558324 114254 558348 114526
rect 558620 114254 558644 114526
rect 558324 8009 558644 114254
rect 561870 116606 562190 219970
rect 561870 116334 561894 116606
rect 562166 116334 562190 116606
rect 558300 7985 558668 8009
rect 558300 7665 558324 7985
rect 558644 7665 558668 7985
rect 558300 7641 558668 7665
rect 554754 6265 555122 6289
rect 554754 5945 554778 6265
rect 555098 5945 555122 6265
rect 561870 6209 562190 116334
rect 565416 119366 565736 222830
rect 565416 119094 565440 119366
rect 565712 119094 565736 119366
rect 565416 6439 565736 119094
rect 568962 121606 569282 225690
rect 568962 121334 568986 121606
rect 569258 121334 569282 121606
rect 565392 6415 565760 6439
rect 568962 6419 569282 121334
rect 572508 124596 572828 229120
rect 576054 226910 576374 234250
rect 573940 226590 576374 226910
rect 572508 124324 572532 124596
rect 572804 124324 572828 124596
rect 572508 6689 572828 124324
rect 576054 131016 576374 226590
rect 576054 130744 576078 131016
rect 576350 130744 576374 131016
rect 576054 9869 576374 130744
rect 576030 9845 576398 9869
rect 576030 9525 576054 9845
rect 576374 9525 576398 9845
rect 576030 9501 576398 9525
rect 572484 6665 572852 6689
rect 554754 5921 555122 5945
rect 561846 6185 562214 6209
rect 561846 5865 561870 6185
rect 562190 5865 562214 6185
rect 565392 6095 565416 6415
rect 565736 6095 565760 6415
rect 565392 6071 565760 6095
rect 568938 6395 569306 6419
rect 568938 6075 568962 6395
rect 569282 6075 569306 6395
rect 572484 6345 572508 6665
rect 572828 6345 572852 6665
rect 572484 6321 572852 6345
rect 568938 6051 569306 6075
rect 561846 5841 562214 5865
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use 8bit_sens  8bit_sens_0
timestamp 1661898952
transform 1 0 52880 0 1 199490
box -110 -750 2810 3340
use adc  adc_0
timestamp 1662180122
transform 1 0 52980 0 1 205530
box 450 -2480 2630 -665
use bias_cell  bias_cell_0
timestamp 1661984010
transform 1 0 24660 0 1 691160
box 790 -2240 11230 -60
use small_array  small_array_0
timestamp 1662181890
transform 1 0 178006 0 1 98263
box 0 -10490 15660 4530
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
rlabel metal1 182035 88193 182035 88193 1 small_array_0/bottom_left_pixel_0/bottom_pixel_0/8bit_sens_0/GND
port 19 n
rlabel metal1 183035 88193 183035 88193 1 small_array_0/bottom_left_pixel_0/bottom_pixel_0/8bit_sens_0/GND
port 19 n
rlabel metal1 185035 88193 185035 88193 1 small_array_0/bottom_left_pixel_0/bottom_pixel_0/8bit_sens_0/GND
port 19 n
rlabel metal1 186035 88193 186035 88193 1 small_array_0/bottom_left_pixel_0/bottom_pixel_0/8bit_sens_0/GND
port 19 n
rlabel metal1 188035 88193 188035 88193 1 small_array_0/bottom_left_pixel_0/bottom_pixel_0/8bit_sens_0/GND
port 19 n
rlabel metal1 189035 88193 189035 88193 1 small_array_0/bottom_left_pixel_0/bottom_pixel_0/8bit_sens_0/GND
port 19 n
rlabel metal1 190035 88193 190035 88193 1 small_array_0/bottom_left_pixel_0/bottom_pixel_0/8bit_sens_0/GND
port 19 n
rlabel metal1 187035 88193 187035 88193 1 small_array_0/bottom_left_pixel_0/bottom_pixel_0/8bit_sens_0/GND
port 19 n
rlabel metal1 184035 88193 184035 88193 1 small_array_0/bottom_left_pixel_0/bottom_pixel_0/8bit_sens_0/GND
port 19 n
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
