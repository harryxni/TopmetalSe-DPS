magic
tech sky130B
magscale 1 2
timestamp 1607731921
<< nwell >>
rect -4172 -1537 4172 1537
<< pmos >>
rect -3976 118 -3856 1318
rect -3798 118 -3678 1318
rect -3620 118 -3500 1318
rect -3442 118 -3322 1318
rect -3264 118 -3144 1318
rect -3086 118 -2966 1318
rect -2908 118 -2788 1318
rect -2730 118 -2610 1318
rect -2552 118 -2432 1318
rect -2374 118 -2254 1318
rect -2196 118 -2076 1318
rect -2018 118 -1898 1318
rect -1840 118 -1720 1318
rect -1662 118 -1542 1318
rect -1484 118 -1364 1318
rect -1306 118 -1186 1318
rect -1128 118 -1008 1318
rect -950 118 -830 1318
rect -772 118 -652 1318
rect -594 118 -474 1318
rect -416 118 -296 1318
rect -238 118 -118 1318
rect -60 118 60 1318
rect 118 118 238 1318
rect 296 118 416 1318
rect 474 118 594 1318
rect 652 118 772 1318
rect 830 118 950 1318
rect 1008 118 1128 1318
rect 1186 118 1306 1318
rect 1364 118 1484 1318
rect 1542 118 1662 1318
rect 1720 118 1840 1318
rect 1898 118 2018 1318
rect 2076 118 2196 1318
rect 2254 118 2374 1318
rect 2432 118 2552 1318
rect 2610 118 2730 1318
rect 2788 118 2908 1318
rect 2966 118 3086 1318
rect 3144 118 3264 1318
rect 3322 118 3442 1318
rect 3500 118 3620 1318
rect 3678 118 3798 1318
rect 3856 118 3976 1318
rect -3976 -1318 -3856 -118
rect -3798 -1318 -3678 -118
rect -3620 -1318 -3500 -118
rect -3442 -1318 -3322 -118
rect -3264 -1318 -3144 -118
rect -3086 -1318 -2966 -118
rect -2908 -1318 -2788 -118
rect -2730 -1318 -2610 -118
rect -2552 -1318 -2432 -118
rect -2374 -1318 -2254 -118
rect -2196 -1318 -2076 -118
rect -2018 -1318 -1898 -118
rect -1840 -1318 -1720 -118
rect -1662 -1318 -1542 -118
rect -1484 -1318 -1364 -118
rect -1306 -1318 -1186 -118
rect -1128 -1318 -1008 -118
rect -950 -1318 -830 -118
rect -772 -1318 -652 -118
rect -594 -1318 -474 -118
rect -416 -1318 -296 -118
rect -238 -1318 -118 -118
rect -60 -1318 60 -118
rect 118 -1318 238 -118
rect 296 -1318 416 -118
rect 474 -1318 594 -118
rect 652 -1318 772 -118
rect 830 -1318 950 -118
rect 1008 -1318 1128 -118
rect 1186 -1318 1306 -118
rect 1364 -1318 1484 -118
rect 1542 -1318 1662 -118
rect 1720 -1318 1840 -118
rect 1898 -1318 2018 -118
rect 2076 -1318 2196 -118
rect 2254 -1318 2374 -118
rect 2432 -1318 2552 -118
rect 2610 -1318 2730 -118
rect 2788 -1318 2908 -118
rect 2966 -1318 3086 -118
rect 3144 -1318 3264 -118
rect 3322 -1318 3442 -118
rect 3500 -1318 3620 -118
rect 3678 -1318 3798 -118
rect 3856 -1318 3976 -118
<< pdiff >>
rect -4034 1306 -3976 1318
rect -4034 130 -4022 1306
rect -3988 130 -3976 1306
rect -4034 118 -3976 130
rect -3856 1306 -3798 1318
rect -3856 130 -3844 1306
rect -3810 130 -3798 1306
rect -3856 118 -3798 130
rect -3678 1306 -3620 1318
rect -3678 130 -3666 1306
rect -3632 130 -3620 1306
rect -3678 118 -3620 130
rect -3500 1306 -3442 1318
rect -3500 130 -3488 1306
rect -3454 130 -3442 1306
rect -3500 118 -3442 130
rect -3322 1306 -3264 1318
rect -3322 130 -3310 1306
rect -3276 130 -3264 1306
rect -3322 118 -3264 130
rect -3144 1306 -3086 1318
rect -3144 130 -3132 1306
rect -3098 130 -3086 1306
rect -3144 118 -3086 130
rect -2966 1306 -2908 1318
rect -2966 130 -2954 1306
rect -2920 130 -2908 1306
rect -2966 118 -2908 130
rect -2788 1306 -2730 1318
rect -2788 130 -2776 1306
rect -2742 130 -2730 1306
rect -2788 118 -2730 130
rect -2610 1306 -2552 1318
rect -2610 130 -2598 1306
rect -2564 130 -2552 1306
rect -2610 118 -2552 130
rect -2432 1306 -2374 1318
rect -2432 130 -2420 1306
rect -2386 130 -2374 1306
rect -2432 118 -2374 130
rect -2254 1306 -2196 1318
rect -2254 130 -2242 1306
rect -2208 130 -2196 1306
rect -2254 118 -2196 130
rect -2076 1306 -2018 1318
rect -2076 130 -2064 1306
rect -2030 130 -2018 1306
rect -2076 118 -2018 130
rect -1898 1306 -1840 1318
rect -1898 130 -1886 1306
rect -1852 130 -1840 1306
rect -1898 118 -1840 130
rect -1720 1306 -1662 1318
rect -1720 130 -1708 1306
rect -1674 130 -1662 1306
rect -1720 118 -1662 130
rect -1542 1306 -1484 1318
rect -1542 130 -1530 1306
rect -1496 130 -1484 1306
rect -1542 118 -1484 130
rect -1364 1306 -1306 1318
rect -1364 130 -1352 1306
rect -1318 130 -1306 1306
rect -1364 118 -1306 130
rect -1186 1306 -1128 1318
rect -1186 130 -1174 1306
rect -1140 130 -1128 1306
rect -1186 118 -1128 130
rect -1008 1306 -950 1318
rect -1008 130 -996 1306
rect -962 130 -950 1306
rect -1008 118 -950 130
rect -830 1306 -772 1318
rect -830 130 -818 1306
rect -784 130 -772 1306
rect -830 118 -772 130
rect -652 1306 -594 1318
rect -652 130 -640 1306
rect -606 130 -594 1306
rect -652 118 -594 130
rect -474 1306 -416 1318
rect -474 130 -462 1306
rect -428 130 -416 1306
rect -474 118 -416 130
rect -296 1306 -238 1318
rect -296 130 -284 1306
rect -250 130 -238 1306
rect -296 118 -238 130
rect -118 1306 -60 1318
rect -118 130 -106 1306
rect -72 130 -60 1306
rect -118 118 -60 130
rect 60 1306 118 1318
rect 60 130 72 1306
rect 106 130 118 1306
rect 60 118 118 130
rect 238 1306 296 1318
rect 238 130 250 1306
rect 284 130 296 1306
rect 238 118 296 130
rect 416 1306 474 1318
rect 416 130 428 1306
rect 462 130 474 1306
rect 416 118 474 130
rect 594 1306 652 1318
rect 594 130 606 1306
rect 640 130 652 1306
rect 594 118 652 130
rect 772 1306 830 1318
rect 772 130 784 1306
rect 818 130 830 1306
rect 772 118 830 130
rect 950 1306 1008 1318
rect 950 130 962 1306
rect 996 130 1008 1306
rect 950 118 1008 130
rect 1128 1306 1186 1318
rect 1128 130 1140 1306
rect 1174 130 1186 1306
rect 1128 118 1186 130
rect 1306 1306 1364 1318
rect 1306 130 1318 1306
rect 1352 130 1364 1306
rect 1306 118 1364 130
rect 1484 1306 1542 1318
rect 1484 130 1496 1306
rect 1530 130 1542 1306
rect 1484 118 1542 130
rect 1662 1306 1720 1318
rect 1662 130 1674 1306
rect 1708 130 1720 1306
rect 1662 118 1720 130
rect 1840 1306 1898 1318
rect 1840 130 1852 1306
rect 1886 130 1898 1306
rect 1840 118 1898 130
rect 2018 1306 2076 1318
rect 2018 130 2030 1306
rect 2064 130 2076 1306
rect 2018 118 2076 130
rect 2196 1306 2254 1318
rect 2196 130 2208 1306
rect 2242 130 2254 1306
rect 2196 118 2254 130
rect 2374 1306 2432 1318
rect 2374 130 2386 1306
rect 2420 130 2432 1306
rect 2374 118 2432 130
rect 2552 1306 2610 1318
rect 2552 130 2564 1306
rect 2598 130 2610 1306
rect 2552 118 2610 130
rect 2730 1306 2788 1318
rect 2730 130 2742 1306
rect 2776 130 2788 1306
rect 2730 118 2788 130
rect 2908 1306 2966 1318
rect 2908 130 2920 1306
rect 2954 130 2966 1306
rect 2908 118 2966 130
rect 3086 1306 3144 1318
rect 3086 130 3098 1306
rect 3132 130 3144 1306
rect 3086 118 3144 130
rect 3264 1306 3322 1318
rect 3264 130 3276 1306
rect 3310 130 3322 1306
rect 3264 118 3322 130
rect 3442 1306 3500 1318
rect 3442 130 3454 1306
rect 3488 130 3500 1306
rect 3442 118 3500 130
rect 3620 1306 3678 1318
rect 3620 130 3632 1306
rect 3666 130 3678 1306
rect 3620 118 3678 130
rect 3798 1306 3856 1318
rect 3798 130 3810 1306
rect 3844 130 3856 1306
rect 3798 118 3856 130
rect 3976 1306 4034 1318
rect 3976 130 3988 1306
rect 4022 130 4034 1306
rect 3976 118 4034 130
rect -4034 -130 -3976 -118
rect -4034 -1306 -4022 -130
rect -3988 -1306 -3976 -130
rect -4034 -1318 -3976 -1306
rect -3856 -130 -3798 -118
rect -3856 -1306 -3844 -130
rect -3810 -1306 -3798 -130
rect -3856 -1318 -3798 -1306
rect -3678 -130 -3620 -118
rect -3678 -1306 -3666 -130
rect -3632 -1306 -3620 -130
rect -3678 -1318 -3620 -1306
rect -3500 -130 -3442 -118
rect -3500 -1306 -3488 -130
rect -3454 -1306 -3442 -130
rect -3500 -1318 -3442 -1306
rect -3322 -130 -3264 -118
rect -3322 -1306 -3310 -130
rect -3276 -1306 -3264 -130
rect -3322 -1318 -3264 -1306
rect -3144 -130 -3086 -118
rect -3144 -1306 -3132 -130
rect -3098 -1306 -3086 -130
rect -3144 -1318 -3086 -1306
rect -2966 -130 -2908 -118
rect -2966 -1306 -2954 -130
rect -2920 -1306 -2908 -130
rect -2966 -1318 -2908 -1306
rect -2788 -130 -2730 -118
rect -2788 -1306 -2776 -130
rect -2742 -1306 -2730 -130
rect -2788 -1318 -2730 -1306
rect -2610 -130 -2552 -118
rect -2610 -1306 -2598 -130
rect -2564 -1306 -2552 -130
rect -2610 -1318 -2552 -1306
rect -2432 -130 -2374 -118
rect -2432 -1306 -2420 -130
rect -2386 -1306 -2374 -130
rect -2432 -1318 -2374 -1306
rect -2254 -130 -2196 -118
rect -2254 -1306 -2242 -130
rect -2208 -1306 -2196 -130
rect -2254 -1318 -2196 -1306
rect -2076 -130 -2018 -118
rect -2076 -1306 -2064 -130
rect -2030 -1306 -2018 -130
rect -2076 -1318 -2018 -1306
rect -1898 -130 -1840 -118
rect -1898 -1306 -1886 -130
rect -1852 -1306 -1840 -130
rect -1898 -1318 -1840 -1306
rect -1720 -130 -1662 -118
rect -1720 -1306 -1708 -130
rect -1674 -1306 -1662 -130
rect -1720 -1318 -1662 -1306
rect -1542 -130 -1484 -118
rect -1542 -1306 -1530 -130
rect -1496 -1306 -1484 -130
rect -1542 -1318 -1484 -1306
rect -1364 -130 -1306 -118
rect -1364 -1306 -1352 -130
rect -1318 -1306 -1306 -130
rect -1364 -1318 -1306 -1306
rect -1186 -130 -1128 -118
rect -1186 -1306 -1174 -130
rect -1140 -1306 -1128 -130
rect -1186 -1318 -1128 -1306
rect -1008 -130 -950 -118
rect -1008 -1306 -996 -130
rect -962 -1306 -950 -130
rect -1008 -1318 -950 -1306
rect -830 -130 -772 -118
rect -830 -1306 -818 -130
rect -784 -1306 -772 -130
rect -830 -1318 -772 -1306
rect -652 -130 -594 -118
rect -652 -1306 -640 -130
rect -606 -1306 -594 -130
rect -652 -1318 -594 -1306
rect -474 -130 -416 -118
rect -474 -1306 -462 -130
rect -428 -1306 -416 -130
rect -474 -1318 -416 -1306
rect -296 -130 -238 -118
rect -296 -1306 -284 -130
rect -250 -1306 -238 -130
rect -296 -1318 -238 -1306
rect -118 -130 -60 -118
rect -118 -1306 -106 -130
rect -72 -1306 -60 -130
rect -118 -1318 -60 -1306
rect 60 -130 118 -118
rect 60 -1306 72 -130
rect 106 -1306 118 -130
rect 60 -1318 118 -1306
rect 238 -130 296 -118
rect 238 -1306 250 -130
rect 284 -1306 296 -130
rect 238 -1318 296 -1306
rect 416 -130 474 -118
rect 416 -1306 428 -130
rect 462 -1306 474 -130
rect 416 -1318 474 -1306
rect 594 -130 652 -118
rect 594 -1306 606 -130
rect 640 -1306 652 -130
rect 594 -1318 652 -1306
rect 772 -130 830 -118
rect 772 -1306 784 -130
rect 818 -1306 830 -130
rect 772 -1318 830 -1306
rect 950 -130 1008 -118
rect 950 -1306 962 -130
rect 996 -1306 1008 -130
rect 950 -1318 1008 -1306
rect 1128 -130 1186 -118
rect 1128 -1306 1140 -130
rect 1174 -1306 1186 -130
rect 1128 -1318 1186 -1306
rect 1306 -130 1364 -118
rect 1306 -1306 1318 -130
rect 1352 -1306 1364 -130
rect 1306 -1318 1364 -1306
rect 1484 -130 1542 -118
rect 1484 -1306 1496 -130
rect 1530 -1306 1542 -130
rect 1484 -1318 1542 -1306
rect 1662 -130 1720 -118
rect 1662 -1306 1674 -130
rect 1708 -1306 1720 -130
rect 1662 -1318 1720 -1306
rect 1840 -130 1898 -118
rect 1840 -1306 1852 -130
rect 1886 -1306 1898 -130
rect 1840 -1318 1898 -1306
rect 2018 -130 2076 -118
rect 2018 -1306 2030 -130
rect 2064 -1306 2076 -130
rect 2018 -1318 2076 -1306
rect 2196 -130 2254 -118
rect 2196 -1306 2208 -130
rect 2242 -1306 2254 -130
rect 2196 -1318 2254 -1306
rect 2374 -130 2432 -118
rect 2374 -1306 2386 -130
rect 2420 -1306 2432 -130
rect 2374 -1318 2432 -1306
rect 2552 -130 2610 -118
rect 2552 -1306 2564 -130
rect 2598 -1306 2610 -130
rect 2552 -1318 2610 -1306
rect 2730 -130 2788 -118
rect 2730 -1306 2742 -130
rect 2776 -1306 2788 -130
rect 2730 -1318 2788 -1306
rect 2908 -130 2966 -118
rect 2908 -1306 2920 -130
rect 2954 -1306 2966 -130
rect 2908 -1318 2966 -1306
rect 3086 -130 3144 -118
rect 3086 -1306 3098 -130
rect 3132 -1306 3144 -130
rect 3086 -1318 3144 -1306
rect 3264 -130 3322 -118
rect 3264 -1306 3276 -130
rect 3310 -1306 3322 -130
rect 3264 -1318 3322 -1306
rect 3442 -130 3500 -118
rect 3442 -1306 3454 -130
rect 3488 -1306 3500 -130
rect 3442 -1318 3500 -1306
rect 3620 -130 3678 -118
rect 3620 -1306 3632 -130
rect 3666 -1306 3678 -130
rect 3620 -1318 3678 -1306
rect 3798 -130 3856 -118
rect 3798 -1306 3810 -130
rect 3844 -1306 3856 -130
rect 3798 -1318 3856 -1306
rect 3976 -130 4034 -118
rect 3976 -1306 3988 -130
rect 4022 -1306 4034 -130
rect 3976 -1318 4034 -1306
<< pdiffc >>
rect -4022 130 -3988 1306
rect -3844 130 -3810 1306
rect -3666 130 -3632 1306
rect -3488 130 -3454 1306
rect -3310 130 -3276 1306
rect -3132 130 -3098 1306
rect -2954 130 -2920 1306
rect -2776 130 -2742 1306
rect -2598 130 -2564 1306
rect -2420 130 -2386 1306
rect -2242 130 -2208 1306
rect -2064 130 -2030 1306
rect -1886 130 -1852 1306
rect -1708 130 -1674 1306
rect -1530 130 -1496 1306
rect -1352 130 -1318 1306
rect -1174 130 -1140 1306
rect -996 130 -962 1306
rect -818 130 -784 1306
rect -640 130 -606 1306
rect -462 130 -428 1306
rect -284 130 -250 1306
rect -106 130 -72 1306
rect 72 130 106 1306
rect 250 130 284 1306
rect 428 130 462 1306
rect 606 130 640 1306
rect 784 130 818 1306
rect 962 130 996 1306
rect 1140 130 1174 1306
rect 1318 130 1352 1306
rect 1496 130 1530 1306
rect 1674 130 1708 1306
rect 1852 130 1886 1306
rect 2030 130 2064 1306
rect 2208 130 2242 1306
rect 2386 130 2420 1306
rect 2564 130 2598 1306
rect 2742 130 2776 1306
rect 2920 130 2954 1306
rect 3098 130 3132 1306
rect 3276 130 3310 1306
rect 3454 130 3488 1306
rect 3632 130 3666 1306
rect 3810 130 3844 1306
rect 3988 130 4022 1306
rect -4022 -1306 -3988 -130
rect -3844 -1306 -3810 -130
rect -3666 -1306 -3632 -130
rect -3488 -1306 -3454 -130
rect -3310 -1306 -3276 -130
rect -3132 -1306 -3098 -130
rect -2954 -1306 -2920 -130
rect -2776 -1306 -2742 -130
rect -2598 -1306 -2564 -130
rect -2420 -1306 -2386 -130
rect -2242 -1306 -2208 -130
rect -2064 -1306 -2030 -130
rect -1886 -1306 -1852 -130
rect -1708 -1306 -1674 -130
rect -1530 -1306 -1496 -130
rect -1352 -1306 -1318 -130
rect -1174 -1306 -1140 -130
rect -996 -1306 -962 -130
rect -818 -1306 -784 -130
rect -640 -1306 -606 -130
rect -462 -1306 -428 -130
rect -284 -1306 -250 -130
rect -106 -1306 -72 -130
rect 72 -1306 106 -130
rect 250 -1306 284 -130
rect 428 -1306 462 -130
rect 606 -1306 640 -130
rect 784 -1306 818 -130
rect 962 -1306 996 -130
rect 1140 -1306 1174 -130
rect 1318 -1306 1352 -130
rect 1496 -1306 1530 -130
rect 1674 -1306 1708 -130
rect 1852 -1306 1886 -130
rect 2030 -1306 2064 -130
rect 2208 -1306 2242 -130
rect 2386 -1306 2420 -130
rect 2564 -1306 2598 -130
rect 2742 -1306 2776 -130
rect 2920 -1306 2954 -130
rect 3098 -1306 3132 -130
rect 3276 -1306 3310 -130
rect 3454 -1306 3488 -130
rect 3632 -1306 3666 -130
rect 3810 -1306 3844 -130
rect 3988 -1306 4022 -130
<< nsubdiff >>
rect -4136 1467 -4040 1501
rect 4040 1467 4136 1501
rect -4136 1405 -4102 1467
rect 4102 1405 4136 1467
rect -4136 -1467 -4102 -1405
rect 4102 -1467 4136 -1405
rect -4136 -1501 -4040 -1467
rect 4040 -1501 4136 -1467
<< nsubdiffcont >>
rect -4040 1467 4040 1501
rect -4136 -1405 -4102 1405
rect 4102 -1405 4136 1405
rect -4040 -1501 4040 -1467
<< poly >>
rect -3976 1399 -3856 1415
rect -3976 1365 -3960 1399
rect -3872 1365 -3856 1399
rect -3976 1318 -3856 1365
rect -3798 1399 -3678 1415
rect -3798 1365 -3782 1399
rect -3694 1365 -3678 1399
rect -3798 1318 -3678 1365
rect -3620 1399 -3500 1415
rect -3620 1365 -3604 1399
rect -3516 1365 -3500 1399
rect -3620 1318 -3500 1365
rect -3442 1399 -3322 1415
rect -3442 1365 -3426 1399
rect -3338 1365 -3322 1399
rect -3442 1318 -3322 1365
rect -3264 1399 -3144 1415
rect -3264 1365 -3248 1399
rect -3160 1365 -3144 1399
rect -3264 1318 -3144 1365
rect -3086 1399 -2966 1415
rect -3086 1365 -3070 1399
rect -2982 1365 -2966 1399
rect -3086 1318 -2966 1365
rect -2908 1399 -2788 1415
rect -2908 1365 -2892 1399
rect -2804 1365 -2788 1399
rect -2908 1318 -2788 1365
rect -2730 1399 -2610 1415
rect -2730 1365 -2714 1399
rect -2626 1365 -2610 1399
rect -2730 1318 -2610 1365
rect -2552 1399 -2432 1415
rect -2552 1365 -2536 1399
rect -2448 1365 -2432 1399
rect -2552 1318 -2432 1365
rect -2374 1399 -2254 1415
rect -2374 1365 -2358 1399
rect -2270 1365 -2254 1399
rect -2374 1318 -2254 1365
rect -2196 1399 -2076 1415
rect -2196 1365 -2180 1399
rect -2092 1365 -2076 1399
rect -2196 1318 -2076 1365
rect -2018 1399 -1898 1415
rect -2018 1365 -2002 1399
rect -1914 1365 -1898 1399
rect -2018 1318 -1898 1365
rect -1840 1399 -1720 1415
rect -1840 1365 -1824 1399
rect -1736 1365 -1720 1399
rect -1840 1318 -1720 1365
rect -1662 1399 -1542 1415
rect -1662 1365 -1646 1399
rect -1558 1365 -1542 1399
rect -1662 1318 -1542 1365
rect -1484 1399 -1364 1415
rect -1484 1365 -1468 1399
rect -1380 1365 -1364 1399
rect -1484 1318 -1364 1365
rect -1306 1399 -1186 1415
rect -1306 1365 -1290 1399
rect -1202 1365 -1186 1399
rect -1306 1318 -1186 1365
rect -1128 1399 -1008 1415
rect -1128 1365 -1112 1399
rect -1024 1365 -1008 1399
rect -1128 1318 -1008 1365
rect -950 1399 -830 1415
rect -950 1365 -934 1399
rect -846 1365 -830 1399
rect -950 1318 -830 1365
rect -772 1399 -652 1415
rect -772 1365 -756 1399
rect -668 1365 -652 1399
rect -772 1318 -652 1365
rect -594 1399 -474 1415
rect -594 1365 -578 1399
rect -490 1365 -474 1399
rect -594 1318 -474 1365
rect -416 1399 -296 1415
rect -416 1365 -400 1399
rect -312 1365 -296 1399
rect -416 1318 -296 1365
rect -238 1399 -118 1415
rect -238 1365 -222 1399
rect -134 1365 -118 1399
rect -238 1318 -118 1365
rect -60 1399 60 1415
rect -60 1365 -44 1399
rect 44 1365 60 1399
rect -60 1318 60 1365
rect 118 1399 238 1415
rect 118 1365 134 1399
rect 222 1365 238 1399
rect 118 1318 238 1365
rect 296 1399 416 1415
rect 296 1365 312 1399
rect 400 1365 416 1399
rect 296 1318 416 1365
rect 474 1399 594 1415
rect 474 1365 490 1399
rect 578 1365 594 1399
rect 474 1318 594 1365
rect 652 1399 772 1415
rect 652 1365 668 1399
rect 756 1365 772 1399
rect 652 1318 772 1365
rect 830 1399 950 1415
rect 830 1365 846 1399
rect 934 1365 950 1399
rect 830 1318 950 1365
rect 1008 1399 1128 1415
rect 1008 1365 1024 1399
rect 1112 1365 1128 1399
rect 1008 1318 1128 1365
rect 1186 1399 1306 1415
rect 1186 1365 1202 1399
rect 1290 1365 1306 1399
rect 1186 1318 1306 1365
rect 1364 1399 1484 1415
rect 1364 1365 1380 1399
rect 1468 1365 1484 1399
rect 1364 1318 1484 1365
rect 1542 1399 1662 1415
rect 1542 1365 1558 1399
rect 1646 1365 1662 1399
rect 1542 1318 1662 1365
rect 1720 1399 1840 1415
rect 1720 1365 1736 1399
rect 1824 1365 1840 1399
rect 1720 1318 1840 1365
rect 1898 1399 2018 1415
rect 1898 1365 1914 1399
rect 2002 1365 2018 1399
rect 1898 1318 2018 1365
rect 2076 1399 2196 1415
rect 2076 1365 2092 1399
rect 2180 1365 2196 1399
rect 2076 1318 2196 1365
rect 2254 1399 2374 1415
rect 2254 1365 2270 1399
rect 2358 1365 2374 1399
rect 2254 1318 2374 1365
rect 2432 1399 2552 1415
rect 2432 1365 2448 1399
rect 2536 1365 2552 1399
rect 2432 1318 2552 1365
rect 2610 1399 2730 1415
rect 2610 1365 2626 1399
rect 2714 1365 2730 1399
rect 2610 1318 2730 1365
rect 2788 1399 2908 1415
rect 2788 1365 2804 1399
rect 2892 1365 2908 1399
rect 2788 1318 2908 1365
rect 2966 1399 3086 1415
rect 2966 1365 2982 1399
rect 3070 1365 3086 1399
rect 2966 1318 3086 1365
rect 3144 1399 3264 1415
rect 3144 1365 3160 1399
rect 3248 1365 3264 1399
rect 3144 1318 3264 1365
rect 3322 1399 3442 1415
rect 3322 1365 3338 1399
rect 3426 1365 3442 1399
rect 3322 1318 3442 1365
rect 3500 1399 3620 1415
rect 3500 1365 3516 1399
rect 3604 1365 3620 1399
rect 3500 1318 3620 1365
rect 3678 1399 3798 1415
rect 3678 1365 3694 1399
rect 3782 1365 3798 1399
rect 3678 1318 3798 1365
rect 3856 1399 3976 1415
rect 3856 1365 3872 1399
rect 3960 1365 3976 1399
rect 3856 1318 3976 1365
rect -3976 71 -3856 118
rect -3976 37 -3960 71
rect -3872 37 -3856 71
rect -3976 21 -3856 37
rect -3798 71 -3678 118
rect -3798 37 -3782 71
rect -3694 37 -3678 71
rect -3798 21 -3678 37
rect -3620 71 -3500 118
rect -3620 37 -3604 71
rect -3516 37 -3500 71
rect -3620 21 -3500 37
rect -3442 71 -3322 118
rect -3442 37 -3426 71
rect -3338 37 -3322 71
rect -3442 21 -3322 37
rect -3264 71 -3144 118
rect -3264 37 -3248 71
rect -3160 37 -3144 71
rect -3264 21 -3144 37
rect -3086 71 -2966 118
rect -3086 37 -3070 71
rect -2982 37 -2966 71
rect -3086 21 -2966 37
rect -2908 71 -2788 118
rect -2908 37 -2892 71
rect -2804 37 -2788 71
rect -2908 21 -2788 37
rect -2730 71 -2610 118
rect -2730 37 -2714 71
rect -2626 37 -2610 71
rect -2730 21 -2610 37
rect -2552 71 -2432 118
rect -2552 37 -2536 71
rect -2448 37 -2432 71
rect -2552 21 -2432 37
rect -2374 71 -2254 118
rect -2374 37 -2358 71
rect -2270 37 -2254 71
rect -2374 21 -2254 37
rect -2196 71 -2076 118
rect -2196 37 -2180 71
rect -2092 37 -2076 71
rect -2196 21 -2076 37
rect -2018 71 -1898 118
rect -2018 37 -2002 71
rect -1914 37 -1898 71
rect -2018 21 -1898 37
rect -1840 71 -1720 118
rect -1840 37 -1824 71
rect -1736 37 -1720 71
rect -1840 21 -1720 37
rect -1662 71 -1542 118
rect -1662 37 -1646 71
rect -1558 37 -1542 71
rect -1662 21 -1542 37
rect -1484 71 -1364 118
rect -1484 37 -1468 71
rect -1380 37 -1364 71
rect -1484 21 -1364 37
rect -1306 71 -1186 118
rect -1306 37 -1290 71
rect -1202 37 -1186 71
rect -1306 21 -1186 37
rect -1128 71 -1008 118
rect -1128 37 -1112 71
rect -1024 37 -1008 71
rect -1128 21 -1008 37
rect -950 71 -830 118
rect -950 37 -934 71
rect -846 37 -830 71
rect -950 21 -830 37
rect -772 71 -652 118
rect -772 37 -756 71
rect -668 37 -652 71
rect -772 21 -652 37
rect -594 71 -474 118
rect -594 37 -578 71
rect -490 37 -474 71
rect -594 21 -474 37
rect -416 71 -296 118
rect -416 37 -400 71
rect -312 37 -296 71
rect -416 21 -296 37
rect -238 71 -118 118
rect -238 37 -222 71
rect -134 37 -118 71
rect -238 21 -118 37
rect -60 71 60 118
rect -60 37 -44 71
rect 44 37 60 71
rect -60 21 60 37
rect 118 71 238 118
rect 118 37 134 71
rect 222 37 238 71
rect 118 21 238 37
rect 296 71 416 118
rect 296 37 312 71
rect 400 37 416 71
rect 296 21 416 37
rect 474 71 594 118
rect 474 37 490 71
rect 578 37 594 71
rect 474 21 594 37
rect 652 71 772 118
rect 652 37 668 71
rect 756 37 772 71
rect 652 21 772 37
rect 830 71 950 118
rect 830 37 846 71
rect 934 37 950 71
rect 830 21 950 37
rect 1008 71 1128 118
rect 1008 37 1024 71
rect 1112 37 1128 71
rect 1008 21 1128 37
rect 1186 71 1306 118
rect 1186 37 1202 71
rect 1290 37 1306 71
rect 1186 21 1306 37
rect 1364 71 1484 118
rect 1364 37 1380 71
rect 1468 37 1484 71
rect 1364 21 1484 37
rect 1542 71 1662 118
rect 1542 37 1558 71
rect 1646 37 1662 71
rect 1542 21 1662 37
rect 1720 71 1840 118
rect 1720 37 1736 71
rect 1824 37 1840 71
rect 1720 21 1840 37
rect 1898 71 2018 118
rect 1898 37 1914 71
rect 2002 37 2018 71
rect 1898 21 2018 37
rect 2076 71 2196 118
rect 2076 37 2092 71
rect 2180 37 2196 71
rect 2076 21 2196 37
rect 2254 71 2374 118
rect 2254 37 2270 71
rect 2358 37 2374 71
rect 2254 21 2374 37
rect 2432 71 2552 118
rect 2432 37 2448 71
rect 2536 37 2552 71
rect 2432 21 2552 37
rect 2610 71 2730 118
rect 2610 37 2626 71
rect 2714 37 2730 71
rect 2610 21 2730 37
rect 2788 71 2908 118
rect 2788 37 2804 71
rect 2892 37 2908 71
rect 2788 21 2908 37
rect 2966 71 3086 118
rect 2966 37 2982 71
rect 3070 37 3086 71
rect 2966 21 3086 37
rect 3144 71 3264 118
rect 3144 37 3160 71
rect 3248 37 3264 71
rect 3144 21 3264 37
rect 3322 71 3442 118
rect 3322 37 3338 71
rect 3426 37 3442 71
rect 3322 21 3442 37
rect 3500 71 3620 118
rect 3500 37 3516 71
rect 3604 37 3620 71
rect 3500 21 3620 37
rect 3678 71 3798 118
rect 3678 37 3694 71
rect 3782 37 3798 71
rect 3678 21 3798 37
rect 3856 71 3976 118
rect 3856 37 3872 71
rect 3960 37 3976 71
rect 3856 21 3976 37
rect -3976 -37 -3856 -21
rect -3976 -71 -3960 -37
rect -3872 -71 -3856 -37
rect -3976 -118 -3856 -71
rect -3798 -37 -3678 -21
rect -3798 -71 -3782 -37
rect -3694 -71 -3678 -37
rect -3798 -118 -3678 -71
rect -3620 -37 -3500 -21
rect -3620 -71 -3604 -37
rect -3516 -71 -3500 -37
rect -3620 -118 -3500 -71
rect -3442 -37 -3322 -21
rect -3442 -71 -3426 -37
rect -3338 -71 -3322 -37
rect -3442 -118 -3322 -71
rect -3264 -37 -3144 -21
rect -3264 -71 -3248 -37
rect -3160 -71 -3144 -37
rect -3264 -118 -3144 -71
rect -3086 -37 -2966 -21
rect -3086 -71 -3070 -37
rect -2982 -71 -2966 -37
rect -3086 -118 -2966 -71
rect -2908 -37 -2788 -21
rect -2908 -71 -2892 -37
rect -2804 -71 -2788 -37
rect -2908 -118 -2788 -71
rect -2730 -37 -2610 -21
rect -2730 -71 -2714 -37
rect -2626 -71 -2610 -37
rect -2730 -118 -2610 -71
rect -2552 -37 -2432 -21
rect -2552 -71 -2536 -37
rect -2448 -71 -2432 -37
rect -2552 -118 -2432 -71
rect -2374 -37 -2254 -21
rect -2374 -71 -2358 -37
rect -2270 -71 -2254 -37
rect -2374 -118 -2254 -71
rect -2196 -37 -2076 -21
rect -2196 -71 -2180 -37
rect -2092 -71 -2076 -37
rect -2196 -118 -2076 -71
rect -2018 -37 -1898 -21
rect -2018 -71 -2002 -37
rect -1914 -71 -1898 -37
rect -2018 -118 -1898 -71
rect -1840 -37 -1720 -21
rect -1840 -71 -1824 -37
rect -1736 -71 -1720 -37
rect -1840 -118 -1720 -71
rect -1662 -37 -1542 -21
rect -1662 -71 -1646 -37
rect -1558 -71 -1542 -37
rect -1662 -118 -1542 -71
rect -1484 -37 -1364 -21
rect -1484 -71 -1468 -37
rect -1380 -71 -1364 -37
rect -1484 -118 -1364 -71
rect -1306 -37 -1186 -21
rect -1306 -71 -1290 -37
rect -1202 -71 -1186 -37
rect -1306 -118 -1186 -71
rect -1128 -37 -1008 -21
rect -1128 -71 -1112 -37
rect -1024 -71 -1008 -37
rect -1128 -118 -1008 -71
rect -950 -37 -830 -21
rect -950 -71 -934 -37
rect -846 -71 -830 -37
rect -950 -118 -830 -71
rect -772 -37 -652 -21
rect -772 -71 -756 -37
rect -668 -71 -652 -37
rect -772 -118 -652 -71
rect -594 -37 -474 -21
rect -594 -71 -578 -37
rect -490 -71 -474 -37
rect -594 -118 -474 -71
rect -416 -37 -296 -21
rect -416 -71 -400 -37
rect -312 -71 -296 -37
rect -416 -118 -296 -71
rect -238 -37 -118 -21
rect -238 -71 -222 -37
rect -134 -71 -118 -37
rect -238 -118 -118 -71
rect -60 -37 60 -21
rect -60 -71 -44 -37
rect 44 -71 60 -37
rect -60 -118 60 -71
rect 118 -37 238 -21
rect 118 -71 134 -37
rect 222 -71 238 -37
rect 118 -118 238 -71
rect 296 -37 416 -21
rect 296 -71 312 -37
rect 400 -71 416 -37
rect 296 -118 416 -71
rect 474 -37 594 -21
rect 474 -71 490 -37
rect 578 -71 594 -37
rect 474 -118 594 -71
rect 652 -37 772 -21
rect 652 -71 668 -37
rect 756 -71 772 -37
rect 652 -118 772 -71
rect 830 -37 950 -21
rect 830 -71 846 -37
rect 934 -71 950 -37
rect 830 -118 950 -71
rect 1008 -37 1128 -21
rect 1008 -71 1024 -37
rect 1112 -71 1128 -37
rect 1008 -118 1128 -71
rect 1186 -37 1306 -21
rect 1186 -71 1202 -37
rect 1290 -71 1306 -37
rect 1186 -118 1306 -71
rect 1364 -37 1484 -21
rect 1364 -71 1380 -37
rect 1468 -71 1484 -37
rect 1364 -118 1484 -71
rect 1542 -37 1662 -21
rect 1542 -71 1558 -37
rect 1646 -71 1662 -37
rect 1542 -118 1662 -71
rect 1720 -37 1840 -21
rect 1720 -71 1736 -37
rect 1824 -71 1840 -37
rect 1720 -118 1840 -71
rect 1898 -37 2018 -21
rect 1898 -71 1914 -37
rect 2002 -71 2018 -37
rect 1898 -118 2018 -71
rect 2076 -37 2196 -21
rect 2076 -71 2092 -37
rect 2180 -71 2196 -37
rect 2076 -118 2196 -71
rect 2254 -37 2374 -21
rect 2254 -71 2270 -37
rect 2358 -71 2374 -37
rect 2254 -118 2374 -71
rect 2432 -37 2552 -21
rect 2432 -71 2448 -37
rect 2536 -71 2552 -37
rect 2432 -118 2552 -71
rect 2610 -37 2730 -21
rect 2610 -71 2626 -37
rect 2714 -71 2730 -37
rect 2610 -118 2730 -71
rect 2788 -37 2908 -21
rect 2788 -71 2804 -37
rect 2892 -71 2908 -37
rect 2788 -118 2908 -71
rect 2966 -37 3086 -21
rect 2966 -71 2982 -37
rect 3070 -71 3086 -37
rect 2966 -118 3086 -71
rect 3144 -37 3264 -21
rect 3144 -71 3160 -37
rect 3248 -71 3264 -37
rect 3144 -118 3264 -71
rect 3322 -37 3442 -21
rect 3322 -71 3338 -37
rect 3426 -71 3442 -37
rect 3322 -118 3442 -71
rect 3500 -37 3620 -21
rect 3500 -71 3516 -37
rect 3604 -71 3620 -37
rect 3500 -118 3620 -71
rect 3678 -37 3798 -21
rect 3678 -71 3694 -37
rect 3782 -71 3798 -37
rect 3678 -118 3798 -71
rect 3856 -37 3976 -21
rect 3856 -71 3872 -37
rect 3960 -71 3976 -37
rect 3856 -118 3976 -71
rect -3976 -1365 -3856 -1318
rect -3976 -1399 -3960 -1365
rect -3872 -1399 -3856 -1365
rect -3976 -1415 -3856 -1399
rect -3798 -1365 -3678 -1318
rect -3798 -1399 -3782 -1365
rect -3694 -1399 -3678 -1365
rect -3798 -1415 -3678 -1399
rect -3620 -1365 -3500 -1318
rect -3620 -1399 -3604 -1365
rect -3516 -1399 -3500 -1365
rect -3620 -1415 -3500 -1399
rect -3442 -1365 -3322 -1318
rect -3442 -1399 -3426 -1365
rect -3338 -1399 -3322 -1365
rect -3442 -1415 -3322 -1399
rect -3264 -1365 -3144 -1318
rect -3264 -1399 -3248 -1365
rect -3160 -1399 -3144 -1365
rect -3264 -1415 -3144 -1399
rect -3086 -1365 -2966 -1318
rect -3086 -1399 -3070 -1365
rect -2982 -1399 -2966 -1365
rect -3086 -1415 -2966 -1399
rect -2908 -1365 -2788 -1318
rect -2908 -1399 -2892 -1365
rect -2804 -1399 -2788 -1365
rect -2908 -1415 -2788 -1399
rect -2730 -1365 -2610 -1318
rect -2730 -1399 -2714 -1365
rect -2626 -1399 -2610 -1365
rect -2730 -1415 -2610 -1399
rect -2552 -1365 -2432 -1318
rect -2552 -1399 -2536 -1365
rect -2448 -1399 -2432 -1365
rect -2552 -1415 -2432 -1399
rect -2374 -1365 -2254 -1318
rect -2374 -1399 -2358 -1365
rect -2270 -1399 -2254 -1365
rect -2374 -1415 -2254 -1399
rect -2196 -1365 -2076 -1318
rect -2196 -1399 -2180 -1365
rect -2092 -1399 -2076 -1365
rect -2196 -1415 -2076 -1399
rect -2018 -1365 -1898 -1318
rect -2018 -1399 -2002 -1365
rect -1914 -1399 -1898 -1365
rect -2018 -1415 -1898 -1399
rect -1840 -1365 -1720 -1318
rect -1840 -1399 -1824 -1365
rect -1736 -1399 -1720 -1365
rect -1840 -1415 -1720 -1399
rect -1662 -1365 -1542 -1318
rect -1662 -1399 -1646 -1365
rect -1558 -1399 -1542 -1365
rect -1662 -1415 -1542 -1399
rect -1484 -1365 -1364 -1318
rect -1484 -1399 -1468 -1365
rect -1380 -1399 -1364 -1365
rect -1484 -1415 -1364 -1399
rect -1306 -1365 -1186 -1318
rect -1306 -1399 -1290 -1365
rect -1202 -1399 -1186 -1365
rect -1306 -1415 -1186 -1399
rect -1128 -1365 -1008 -1318
rect -1128 -1399 -1112 -1365
rect -1024 -1399 -1008 -1365
rect -1128 -1415 -1008 -1399
rect -950 -1365 -830 -1318
rect -950 -1399 -934 -1365
rect -846 -1399 -830 -1365
rect -950 -1415 -830 -1399
rect -772 -1365 -652 -1318
rect -772 -1399 -756 -1365
rect -668 -1399 -652 -1365
rect -772 -1415 -652 -1399
rect -594 -1365 -474 -1318
rect -594 -1399 -578 -1365
rect -490 -1399 -474 -1365
rect -594 -1415 -474 -1399
rect -416 -1365 -296 -1318
rect -416 -1399 -400 -1365
rect -312 -1399 -296 -1365
rect -416 -1415 -296 -1399
rect -238 -1365 -118 -1318
rect -238 -1399 -222 -1365
rect -134 -1399 -118 -1365
rect -238 -1415 -118 -1399
rect -60 -1365 60 -1318
rect -60 -1399 -44 -1365
rect 44 -1399 60 -1365
rect -60 -1415 60 -1399
rect 118 -1365 238 -1318
rect 118 -1399 134 -1365
rect 222 -1399 238 -1365
rect 118 -1415 238 -1399
rect 296 -1365 416 -1318
rect 296 -1399 312 -1365
rect 400 -1399 416 -1365
rect 296 -1415 416 -1399
rect 474 -1365 594 -1318
rect 474 -1399 490 -1365
rect 578 -1399 594 -1365
rect 474 -1415 594 -1399
rect 652 -1365 772 -1318
rect 652 -1399 668 -1365
rect 756 -1399 772 -1365
rect 652 -1415 772 -1399
rect 830 -1365 950 -1318
rect 830 -1399 846 -1365
rect 934 -1399 950 -1365
rect 830 -1415 950 -1399
rect 1008 -1365 1128 -1318
rect 1008 -1399 1024 -1365
rect 1112 -1399 1128 -1365
rect 1008 -1415 1128 -1399
rect 1186 -1365 1306 -1318
rect 1186 -1399 1202 -1365
rect 1290 -1399 1306 -1365
rect 1186 -1415 1306 -1399
rect 1364 -1365 1484 -1318
rect 1364 -1399 1380 -1365
rect 1468 -1399 1484 -1365
rect 1364 -1415 1484 -1399
rect 1542 -1365 1662 -1318
rect 1542 -1399 1558 -1365
rect 1646 -1399 1662 -1365
rect 1542 -1415 1662 -1399
rect 1720 -1365 1840 -1318
rect 1720 -1399 1736 -1365
rect 1824 -1399 1840 -1365
rect 1720 -1415 1840 -1399
rect 1898 -1365 2018 -1318
rect 1898 -1399 1914 -1365
rect 2002 -1399 2018 -1365
rect 1898 -1415 2018 -1399
rect 2076 -1365 2196 -1318
rect 2076 -1399 2092 -1365
rect 2180 -1399 2196 -1365
rect 2076 -1415 2196 -1399
rect 2254 -1365 2374 -1318
rect 2254 -1399 2270 -1365
rect 2358 -1399 2374 -1365
rect 2254 -1415 2374 -1399
rect 2432 -1365 2552 -1318
rect 2432 -1399 2448 -1365
rect 2536 -1399 2552 -1365
rect 2432 -1415 2552 -1399
rect 2610 -1365 2730 -1318
rect 2610 -1399 2626 -1365
rect 2714 -1399 2730 -1365
rect 2610 -1415 2730 -1399
rect 2788 -1365 2908 -1318
rect 2788 -1399 2804 -1365
rect 2892 -1399 2908 -1365
rect 2788 -1415 2908 -1399
rect 2966 -1365 3086 -1318
rect 2966 -1399 2982 -1365
rect 3070 -1399 3086 -1365
rect 2966 -1415 3086 -1399
rect 3144 -1365 3264 -1318
rect 3144 -1399 3160 -1365
rect 3248 -1399 3264 -1365
rect 3144 -1415 3264 -1399
rect 3322 -1365 3442 -1318
rect 3322 -1399 3338 -1365
rect 3426 -1399 3442 -1365
rect 3322 -1415 3442 -1399
rect 3500 -1365 3620 -1318
rect 3500 -1399 3516 -1365
rect 3604 -1399 3620 -1365
rect 3500 -1415 3620 -1399
rect 3678 -1365 3798 -1318
rect 3678 -1399 3694 -1365
rect 3782 -1399 3798 -1365
rect 3678 -1415 3798 -1399
rect 3856 -1365 3976 -1318
rect 3856 -1399 3872 -1365
rect 3960 -1399 3976 -1365
rect 3856 -1415 3976 -1399
<< polycont >>
rect -3960 1365 -3872 1399
rect -3782 1365 -3694 1399
rect -3604 1365 -3516 1399
rect -3426 1365 -3338 1399
rect -3248 1365 -3160 1399
rect -3070 1365 -2982 1399
rect -2892 1365 -2804 1399
rect -2714 1365 -2626 1399
rect -2536 1365 -2448 1399
rect -2358 1365 -2270 1399
rect -2180 1365 -2092 1399
rect -2002 1365 -1914 1399
rect -1824 1365 -1736 1399
rect -1646 1365 -1558 1399
rect -1468 1365 -1380 1399
rect -1290 1365 -1202 1399
rect -1112 1365 -1024 1399
rect -934 1365 -846 1399
rect -756 1365 -668 1399
rect -578 1365 -490 1399
rect -400 1365 -312 1399
rect -222 1365 -134 1399
rect -44 1365 44 1399
rect 134 1365 222 1399
rect 312 1365 400 1399
rect 490 1365 578 1399
rect 668 1365 756 1399
rect 846 1365 934 1399
rect 1024 1365 1112 1399
rect 1202 1365 1290 1399
rect 1380 1365 1468 1399
rect 1558 1365 1646 1399
rect 1736 1365 1824 1399
rect 1914 1365 2002 1399
rect 2092 1365 2180 1399
rect 2270 1365 2358 1399
rect 2448 1365 2536 1399
rect 2626 1365 2714 1399
rect 2804 1365 2892 1399
rect 2982 1365 3070 1399
rect 3160 1365 3248 1399
rect 3338 1365 3426 1399
rect 3516 1365 3604 1399
rect 3694 1365 3782 1399
rect 3872 1365 3960 1399
rect -3960 37 -3872 71
rect -3782 37 -3694 71
rect -3604 37 -3516 71
rect -3426 37 -3338 71
rect -3248 37 -3160 71
rect -3070 37 -2982 71
rect -2892 37 -2804 71
rect -2714 37 -2626 71
rect -2536 37 -2448 71
rect -2358 37 -2270 71
rect -2180 37 -2092 71
rect -2002 37 -1914 71
rect -1824 37 -1736 71
rect -1646 37 -1558 71
rect -1468 37 -1380 71
rect -1290 37 -1202 71
rect -1112 37 -1024 71
rect -934 37 -846 71
rect -756 37 -668 71
rect -578 37 -490 71
rect -400 37 -312 71
rect -222 37 -134 71
rect -44 37 44 71
rect 134 37 222 71
rect 312 37 400 71
rect 490 37 578 71
rect 668 37 756 71
rect 846 37 934 71
rect 1024 37 1112 71
rect 1202 37 1290 71
rect 1380 37 1468 71
rect 1558 37 1646 71
rect 1736 37 1824 71
rect 1914 37 2002 71
rect 2092 37 2180 71
rect 2270 37 2358 71
rect 2448 37 2536 71
rect 2626 37 2714 71
rect 2804 37 2892 71
rect 2982 37 3070 71
rect 3160 37 3248 71
rect 3338 37 3426 71
rect 3516 37 3604 71
rect 3694 37 3782 71
rect 3872 37 3960 71
rect -3960 -71 -3872 -37
rect -3782 -71 -3694 -37
rect -3604 -71 -3516 -37
rect -3426 -71 -3338 -37
rect -3248 -71 -3160 -37
rect -3070 -71 -2982 -37
rect -2892 -71 -2804 -37
rect -2714 -71 -2626 -37
rect -2536 -71 -2448 -37
rect -2358 -71 -2270 -37
rect -2180 -71 -2092 -37
rect -2002 -71 -1914 -37
rect -1824 -71 -1736 -37
rect -1646 -71 -1558 -37
rect -1468 -71 -1380 -37
rect -1290 -71 -1202 -37
rect -1112 -71 -1024 -37
rect -934 -71 -846 -37
rect -756 -71 -668 -37
rect -578 -71 -490 -37
rect -400 -71 -312 -37
rect -222 -71 -134 -37
rect -44 -71 44 -37
rect 134 -71 222 -37
rect 312 -71 400 -37
rect 490 -71 578 -37
rect 668 -71 756 -37
rect 846 -71 934 -37
rect 1024 -71 1112 -37
rect 1202 -71 1290 -37
rect 1380 -71 1468 -37
rect 1558 -71 1646 -37
rect 1736 -71 1824 -37
rect 1914 -71 2002 -37
rect 2092 -71 2180 -37
rect 2270 -71 2358 -37
rect 2448 -71 2536 -37
rect 2626 -71 2714 -37
rect 2804 -71 2892 -37
rect 2982 -71 3070 -37
rect 3160 -71 3248 -37
rect 3338 -71 3426 -37
rect 3516 -71 3604 -37
rect 3694 -71 3782 -37
rect 3872 -71 3960 -37
rect -3960 -1399 -3872 -1365
rect -3782 -1399 -3694 -1365
rect -3604 -1399 -3516 -1365
rect -3426 -1399 -3338 -1365
rect -3248 -1399 -3160 -1365
rect -3070 -1399 -2982 -1365
rect -2892 -1399 -2804 -1365
rect -2714 -1399 -2626 -1365
rect -2536 -1399 -2448 -1365
rect -2358 -1399 -2270 -1365
rect -2180 -1399 -2092 -1365
rect -2002 -1399 -1914 -1365
rect -1824 -1399 -1736 -1365
rect -1646 -1399 -1558 -1365
rect -1468 -1399 -1380 -1365
rect -1290 -1399 -1202 -1365
rect -1112 -1399 -1024 -1365
rect -934 -1399 -846 -1365
rect -756 -1399 -668 -1365
rect -578 -1399 -490 -1365
rect -400 -1399 -312 -1365
rect -222 -1399 -134 -1365
rect -44 -1399 44 -1365
rect 134 -1399 222 -1365
rect 312 -1399 400 -1365
rect 490 -1399 578 -1365
rect 668 -1399 756 -1365
rect 846 -1399 934 -1365
rect 1024 -1399 1112 -1365
rect 1202 -1399 1290 -1365
rect 1380 -1399 1468 -1365
rect 1558 -1399 1646 -1365
rect 1736 -1399 1824 -1365
rect 1914 -1399 2002 -1365
rect 2092 -1399 2180 -1365
rect 2270 -1399 2358 -1365
rect 2448 -1399 2536 -1365
rect 2626 -1399 2714 -1365
rect 2804 -1399 2892 -1365
rect 2982 -1399 3070 -1365
rect 3160 -1399 3248 -1365
rect 3338 -1399 3426 -1365
rect 3516 -1399 3604 -1365
rect 3694 -1399 3782 -1365
rect 3872 -1399 3960 -1365
<< locali >>
rect -4136 1467 -4040 1501
rect 4040 1467 4136 1501
rect -4136 1405 -4102 1467
rect 4102 1405 4136 1467
rect -3976 1365 -3960 1399
rect -3872 1365 -3856 1399
rect -3798 1365 -3782 1399
rect -3694 1365 -3678 1399
rect -3620 1365 -3604 1399
rect -3516 1365 -3500 1399
rect -3442 1365 -3426 1399
rect -3338 1365 -3322 1399
rect -3264 1365 -3248 1399
rect -3160 1365 -3144 1399
rect -3086 1365 -3070 1399
rect -2982 1365 -2966 1399
rect -2908 1365 -2892 1399
rect -2804 1365 -2788 1399
rect -2730 1365 -2714 1399
rect -2626 1365 -2610 1399
rect -2552 1365 -2536 1399
rect -2448 1365 -2432 1399
rect -2374 1365 -2358 1399
rect -2270 1365 -2254 1399
rect -2196 1365 -2180 1399
rect -2092 1365 -2076 1399
rect -2018 1365 -2002 1399
rect -1914 1365 -1898 1399
rect -1840 1365 -1824 1399
rect -1736 1365 -1720 1399
rect -1662 1365 -1646 1399
rect -1558 1365 -1542 1399
rect -1484 1365 -1468 1399
rect -1380 1365 -1364 1399
rect -1306 1365 -1290 1399
rect -1202 1365 -1186 1399
rect -1128 1365 -1112 1399
rect -1024 1365 -1008 1399
rect -950 1365 -934 1399
rect -846 1365 -830 1399
rect -772 1365 -756 1399
rect -668 1365 -652 1399
rect -594 1365 -578 1399
rect -490 1365 -474 1399
rect -416 1365 -400 1399
rect -312 1365 -296 1399
rect -238 1365 -222 1399
rect -134 1365 -118 1399
rect -60 1365 -44 1399
rect 44 1365 60 1399
rect 118 1365 134 1399
rect 222 1365 238 1399
rect 296 1365 312 1399
rect 400 1365 416 1399
rect 474 1365 490 1399
rect 578 1365 594 1399
rect 652 1365 668 1399
rect 756 1365 772 1399
rect 830 1365 846 1399
rect 934 1365 950 1399
rect 1008 1365 1024 1399
rect 1112 1365 1128 1399
rect 1186 1365 1202 1399
rect 1290 1365 1306 1399
rect 1364 1365 1380 1399
rect 1468 1365 1484 1399
rect 1542 1365 1558 1399
rect 1646 1365 1662 1399
rect 1720 1365 1736 1399
rect 1824 1365 1840 1399
rect 1898 1365 1914 1399
rect 2002 1365 2018 1399
rect 2076 1365 2092 1399
rect 2180 1365 2196 1399
rect 2254 1365 2270 1399
rect 2358 1365 2374 1399
rect 2432 1365 2448 1399
rect 2536 1365 2552 1399
rect 2610 1365 2626 1399
rect 2714 1365 2730 1399
rect 2788 1365 2804 1399
rect 2892 1365 2908 1399
rect 2966 1365 2982 1399
rect 3070 1365 3086 1399
rect 3144 1365 3160 1399
rect 3248 1365 3264 1399
rect 3322 1365 3338 1399
rect 3426 1365 3442 1399
rect 3500 1365 3516 1399
rect 3604 1365 3620 1399
rect 3678 1365 3694 1399
rect 3782 1365 3798 1399
rect 3856 1365 3872 1399
rect 3960 1365 3976 1399
rect -4022 1306 -3988 1322
rect -4022 114 -3988 130
rect -3844 1306 -3810 1322
rect -3844 114 -3810 130
rect -3666 1306 -3632 1322
rect -3666 114 -3632 130
rect -3488 1306 -3454 1322
rect -3488 114 -3454 130
rect -3310 1306 -3276 1322
rect -3310 114 -3276 130
rect -3132 1306 -3098 1322
rect -3132 114 -3098 130
rect -2954 1306 -2920 1322
rect -2954 114 -2920 130
rect -2776 1306 -2742 1322
rect -2776 114 -2742 130
rect -2598 1306 -2564 1322
rect -2598 114 -2564 130
rect -2420 1306 -2386 1322
rect -2420 114 -2386 130
rect -2242 1306 -2208 1322
rect -2242 114 -2208 130
rect -2064 1306 -2030 1322
rect -2064 114 -2030 130
rect -1886 1306 -1852 1322
rect -1886 114 -1852 130
rect -1708 1306 -1674 1322
rect -1708 114 -1674 130
rect -1530 1306 -1496 1322
rect -1530 114 -1496 130
rect -1352 1306 -1318 1322
rect -1352 114 -1318 130
rect -1174 1306 -1140 1322
rect -1174 114 -1140 130
rect -996 1306 -962 1322
rect -996 114 -962 130
rect -818 1306 -784 1322
rect -818 114 -784 130
rect -640 1306 -606 1322
rect -640 114 -606 130
rect -462 1306 -428 1322
rect -462 114 -428 130
rect -284 1306 -250 1322
rect -284 114 -250 130
rect -106 1306 -72 1322
rect -106 114 -72 130
rect 72 1306 106 1322
rect 72 114 106 130
rect 250 1306 284 1322
rect 250 114 284 130
rect 428 1306 462 1322
rect 428 114 462 130
rect 606 1306 640 1322
rect 606 114 640 130
rect 784 1306 818 1322
rect 784 114 818 130
rect 962 1306 996 1322
rect 962 114 996 130
rect 1140 1306 1174 1322
rect 1140 114 1174 130
rect 1318 1306 1352 1322
rect 1318 114 1352 130
rect 1496 1306 1530 1322
rect 1496 114 1530 130
rect 1674 1306 1708 1322
rect 1674 114 1708 130
rect 1852 1306 1886 1322
rect 1852 114 1886 130
rect 2030 1306 2064 1322
rect 2030 114 2064 130
rect 2208 1306 2242 1322
rect 2208 114 2242 130
rect 2386 1306 2420 1322
rect 2386 114 2420 130
rect 2564 1306 2598 1322
rect 2564 114 2598 130
rect 2742 1306 2776 1322
rect 2742 114 2776 130
rect 2920 1306 2954 1322
rect 2920 114 2954 130
rect 3098 1306 3132 1322
rect 3098 114 3132 130
rect 3276 1306 3310 1322
rect 3276 114 3310 130
rect 3454 1306 3488 1322
rect 3454 114 3488 130
rect 3632 1306 3666 1322
rect 3632 114 3666 130
rect 3810 1306 3844 1322
rect 3810 114 3844 130
rect 3988 1306 4022 1322
rect 3988 114 4022 130
rect -3976 37 -3960 71
rect -3872 37 -3856 71
rect -3798 37 -3782 71
rect -3694 37 -3678 71
rect -3620 37 -3604 71
rect -3516 37 -3500 71
rect -3442 37 -3426 71
rect -3338 37 -3322 71
rect -3264 37 -3248 71
rect -3160 37 -3144 71
rect -3086 37 -3070 71
rect -2982 37 -2966 71
rect -2908 37 -2892 71
rect -2804 37 -2788 71
rect -2730 37 -2714 71
rect -2626 37 -2610 71
rect -2552 37 -2536 71
rect -2448 37 -2432 71
rect -2374 37 -2358 71
rect -2270 37 -2254 71
rect -2196 37 -2180 71
rect -2092 37 -2076 71
rect -2018 37 -2002 71
rect -1914 37 -1898 71
rect -1840 37 -1824 71
rect -1736 37 -1720 71
rect -1662 37 -1646 71
rect -1558 37 -1542 71
rect -1484 37 -1468 71
rect -1380 37 -1364 71
rect -1306 37 -1290 71
rect -1202 37 -1186 71
rect -1128 37 -1112 71
rect -1024 37 -1008 71
rect -950 37 -934 71
rect -846 37 -830 71
rect -772 37 -756 71
rect -668 37 -652 71
rect -594 37 -578 71
rect -490 37 -474 71
rect -416 37 -400 71
rect -312 37 -296 71
rect -238 37 -222 71
rect -134 37 -118 71
rect -60 37 -44 71
rect 44 37 60 71
rect 118 37 134 71
rect 222 37 238 71
rect 296 37 312 71
rect 400 37 416 71
rect 474 37 490 71
rect 578 37 594 71
rect 652 37 668 71
rect 756 37 772 71
rect 830 37 846 71
rect 934 37 950 71
rect 1008 37 1024 71
rect 1112 37 1128 71
rect 1186 37 1202 71
rect 1290 37 1306 71
rect 1364 37 1380 71
rect 1468 37 1484 71
rect 1542 37 1558 71
rect 1646 37 1662 71
rect 1720 37 1736 71
rect 1824 37 1840 71
rect 1898 37 1914 71
rect 2002 37 2018 71
rect 2076 37 2092 71
rect 2180 37 2196 71
rect 2254 37 2270 71
rect 2358 37 2374 71
rect 2432 37 2448 71
rect 2536 37 2552 71
rect 2610 37 2626 71
rect 2714 37 2730 71
rect 2788 37 2804 71
rect 2892 37 2908 71
rect 2966 37 2982 71
rect 3070 37 3086 71
rect 3144 37 3160 71
rect 3248 37 3264 71
rect 3322 37 3338 71
rect 3426 37 3442 71
rect 3500 37 3516 71
rect 3604 37 3620 71
rect 3678 37 3694 71
rect 3782 37 3798 71
rect 3856 37 3872 71
rect 3960 37 3976 71
rect -3976 -71 -3960 -37
rect -3872 -71 -3856 -37
rect -3798 -71 -3782 -37
rect -3694 -71 -3678 -37
rect -3620 -71 -3604 -37
rect -3516 -71 -3500 -37
rect -3442 -71 -3426 -37
rect -3338 -71 -3322 -37
rect -3264 -71 -3248 -37
rect -3160 -71 -3144 -37
rect -3086 -71 -3070 -37
rect -2982 -71 -2966 -37
rect -2908 -71 -2892 -37
rect -2804 -71 -2788 -37
rect -2730 -71 -2714 -37
rect -2626 -71 -2610 -37
rect -2552 -71 -2536 -37
rect -2448 -71 -2432 -37
rect -2374 -71 -2358 -37
rect -2270 -71 -2254 -37
rect -2196 -71 -2180 -37
rect -2092 -71 -2076 -37
rect -2018 -71 -2002 -37
rect -1914 -71 -1898 -37
rect -1840 -71 -1824 -37
rect -1736 -71 -1720 -37
rect -1662 -71 -1646 -37
rect -1558 -71 -1542 -37
rect -1484 -71 -1468 -37
rect -1380 -71 -1364 -37
rect -1306 -71 -1290 -37
rect -1202 -71 -1186 -37
rect -1128 -71 -1112 -37
rect -1024 -71 -1008 -37
rect -950 -71 -934 -37
rect -846 -71 -830 -37
rect -772 -71 -756 -37
rect -668 -71 -652 -37
rect -594 -71 -578 -37
rect -490 -71 -474 -37
rect -416 -71 -400 -37
rect -312 -71 -296 -37
rect -238 -71 -222 -37
rect -134 -71 -118 -37
rect -60 -71 -44 -37
rect 44 -71 60 -37
rect 118 -71 134 -37
rect 222 -71 238 -37
rect 296 -71 312 -37
rect 400 -71 416 -37
rect 474 -71 490 -37
rect 578 -71 594 -37
rect 652 -71 668 -37
rect 756 -71 772 -37
rect 830 -71 846 -37
rect 934 -71 950 -37
rect 1008 -71 1024 -37
rect 1112 -71 1128 -37
rect 1186 -71 1202 -37
rect 1290 -71 1306 -37
rect 1364 -71 1380 -37
rect 1468 -71 1484 -37
rect 1542 -71 1558 -37
rect 1646 -71 1662 -37
rect 1720 -71 1736 -37
rect 1824 -71 1840 -37
rect 1898 -71 1914 -37
rect 2002 -71 2018 -37
rect 2076 -71 2092 -37
rect 2180 -71 2196 -37
rect 2254 -71 2270 -37
rect 2358 -71 2374 -37
rect 2432 -71 2448 -37
rect 2536 -71 2552 -37
rect 2610 -71 2626 -37
rect 2714 -71 2730 -37
rect 2788 -71 2804 -37
rect 2892 -71 2908 -37
rect 2966 -71 2982 -37
rect 3070 -71 3086 -37
rect 3144 -71 3160 -37
rect 3248 -71 3264 -37
rect 3322 -71 3338 -37
rect 3426 -71 3442 -37
rect 3500 -71 3516 -37
rect 3604 -71 3620 -37
rect 3678 -71 3694 -37
rect 3782 -71 3798 -37
rect 3856 -71 3872 -37
rect 3960 -71 3976 -37
rect -4022 -130 -3988 -114
rect -4022 -1322 -3988 -1306
rect -3844 -130 -3810 -114
rect -3844 -1322 -3810 -1306
rect -3666 -130 -3632 -114
rect -3666 -1322 -3632 -1306
rect -3488 -130 -3454 -114
rect -3488 -1322 -3454 -1306
rect -3310 -130 -3276 -114
rect -3310 -1322 -3276 -1306
rect -3132 -130 -3098 -114
rect -3132 -1322 -3098 -1306
rect -2954 -130 -2920 -114
rect -2954 -1322 -2920 -1306
rect -2776 -130 -2742 -114
rect -2776 -1322 -2742 -1306
rect -2598 -130 -2564 -114
rect -2598 -1322 -2564 -1306
rect -2420 -130 -2386 -114
rect -2420 -1322 -2386 -1306
rect -2242 -130 -2208 -114
rect -2242 -1322 -2208 -1306
rect -2064 -130 -2030 -114
rect -2064 -1322 -2030 -1306
rect -1886 -130 -1852 -114
rect -1886 -1322 -1852 -1306
rect -1708 -130 -1674 -114
rect -1708 -1322 -1674 -1306
rect -1530 -130 -1496 -114
rect -1530 -1322 -1496 -1306
rect -1352 -130 -1318 -114
rect -1352 -1322 -1318 -1306
rect -1174 -130 -1140 -114
rect -1174 -1322 -1140 -1306
rect -996 -130 -962 -114
rect -996 -1322 -962 -1306
rect -818 -130 -784 -114
rect -818 -1322 -784 -1306
rect -640 -130 -606 -114
rect -640 -1322 -606 -1306
rect -462 -130 -428 -114
rect -462 -1322 -428 -1306
rect -284 -130 -250 -114
rect -284 -1322 -250 -1306
rect -106 -130 -72 -114
rect -106 -1322 -72 -1306
rect 72 -130 106 -114
rect 72 -1322 106 -1306
rect 250 -130 284 -114
rect 250 -1322 284 -1306
rect 428 -130 462 -114
rect 428 -1322 462 -1306
rect 606 -130 640 -114
rect 606 -1322 640 -1306
rect 784 -130 818 -114
rect 784 -1322 818 -1306
rect 962 -130 996 -114
rect 962 -1322 996 -1306
rect 1140 -130 1174 -114
rect 1140 -1322 1174 -1306
rect 1318 -130 1352 -114
rect 1318 -1322 1352 -1306
rect 1496 -130 1530 -114
rect 1496 -1322 1530 -1306
rect 1674 -130 1708 -114
rect 1674 -1322 1708 -1306
rect 1852 -130 1886 -114
rect 1852 -1322 1886 -1306
rect 2030 -130 2064 -114
rect 2030 -1322 2064 -1306
rect 2208 -130 2242 -114
rect 2208 -1322 2242 -1306
rect 2386 -130 2420 -114
rect 2386 -1322 2420 -1306
rect 2564 -130 2598 -114
rect 2564 -1322 2598 -1306
rect 2742 -130 2776 -114
rect 2742 -1322 2776 -1306
rect 2920 -130 2954 -114
rect 2920 -1322 2954 -1306
rect 3098 -130 3132 -114
rect 3098 -1322 3132 -1306
rect 3276 -130 3310 -114
rect 3276 -1322 3310 -1306
rect 3454 -130 3488 -114
rect 3454 -1322 3488 -1306
rect 3632 -130 3666 -114
rect 3632 -1322 3666 -1306
rect 3810 -130 3844 -114
rect 3810 -1322 3844 -1306
rect 3988 -130 4022 -114
rect 3988 -1322 4022 -1306
rect -3976 -1399 -3960 -1365
rect -3872 -1399 -3856 -1365
rect -3798 -1399 -3782 -1365
rect -3694 -1399 -3678 -1365
rect -3620 -1399 -3604 -1365
rect -3516 -1399 -3500 -1365
rect -3442 -1399 -3426 -1365
rect -3338 -1399 -3322 -1365
rect -3264 -1399 -3248 -1365
rect -3160 -1399 -3144 -1365
rect -3086 -1399 -3070 -1365
rect -2982 -1399 -2966 -1365
rect -2908 -1399 -2892 -1365
rect -2804 -1399 -2788 -1365
rect -2730 -1399 -2714 -1365
rect -2626 -1399 -2610 -1365
rect -2552 -1399 -2536 -1365
rect -2448 -1399 -2432 -1365
rect -2374 -1399 -2358 -1365
rect -2270 -1399 -2254 -1365
rect -2196 -1399 -2180 -1365
rect -2092 -1399 -2076 -1365
rect -2018 -1399 -2002 -1365
rect -1914 -1399 -1898 -1365
rect -1840 -1399 -1824 -1365
rect -1736 -1399 -1720 -1365
rect -1662 -1399 -1646 -1365
rect -1558 -1399 -1542 -1365
rect -1484 -1399 -1468 -1365
rect -1380 -1399 -1364 -1365
rect -1306 -1399 -1290 -1365
rect -1202 -1399 -1186 -1365
rect -1128 -1399 -1112 -1365
rect -1024 -1399 -1008 -1365
rect -950 -1399 -934 -1365
rect -846 -1399 -830 -1365
rect -772 -1399 -756 -1365
rect -668 -1399 -652 -1365
rect -594 -1399 -578 -1365
rect -490 -1399 -474 -1365
rect -416 -1399 -400 -1365
rect -312 -1399 -296 -1365
rect -238 -1399 -222 -1365
rect -134 -1399 -118 -1365
rect -60 -1399 -44 -1365
rect 44 -1399 60 -1365
rect 118 -1399 134 -1365
rect 222 -1399 238 -1365
rect 296 -1399 312 -1365
rect 400 -1399 416 -1365
rect 474 -1399 490 -1365
rect 578 -1399 594 -1365
rect 652 -1399 668 -1365
rect 756 -1399 772 -1365
rect 830 -1399 846 -1365
rect 934 -1399 950 -1365
rect 1008 -1399 1024 -1365
rect 1112 -1399 1128 -1365
rect 1186 -1399 1202 -1365
rect 1290 -1399 1306 -1365
rect 1364 -1399 1380 -1365
rect 1468 -1399 1484 -1365
rect 1542 -1399 1558 -1365
rect 1646 -1399 1662 -1365
rect 1720 -1399 1736 -1365
rect 1824 -1399 1840 -1365
rect 1898 -1399 1914 -1365
rect 2002 -1399 2018 -1365
rect 2076 -1399 2092 -1365
rect 2180 -1399 2196 -1365
rect 2254 -1399 2270 -1365
rect 2358 -1399 2374 -1365
rect 2432 -1399 2448 -1365
rect 2536 -1399 2552 -1365
rect 2610 -1399 2626 -1365
rect 2714 -1399 2730 -1365
rect 2788 -1399 2804 -1365
rect 2892 -1399 2908 -1365
rect 2966 -1399 2982 -1365
rect 3070 -1399 3086 -1365
rect 3144 -1399 3160 -1365
rect 3248 -1399 3264 -1365
rect 3322 -1399 3338 -1365
rect 3426 -1399 3442 -1365
rect 3500 -1399 3516 -1365
rect 3604 -1399 3620 -1365
rect 3678 -1399 3694 -1365
rect 3782 -1399 3798 -1365
rect 3856 -1399 3872 -1365
rect 3960 -1399 3976 -1365
rect -4136 -1467 -4102 -1405
rect 4102 -1467 4136 -1405
rect -4136 -1501 -4040 -1467
rect 4040 -1501 4136 -1467
<< viali >>
rect -3960 1365 -3872 1399
rect -3782 1365 -3694 1399
rect -3604 1365 -3516 1399
rect -3426 1365 -3338 1399
rect -3248 1365 -3160 1399
rect -3070 1365 -2982 1399
rect -2892 1365 -2804 1399
rect -2714 1365 -2626 1399
rect -2536 1365 -2448 1399
rect -2358 1365 -2270 1399
rect -2180 1365 -2092 1399
rect -2002 1365 -1914 1399
rect -1824 1365 -1736 1399
rect -1646 1365 -1558 1399
rect -1468 1365 -1380 1399
rect -1290 1365 -1202 1399
rect -1112 1365 -1024 1399
rect -934 1365 -846 1399
rect -756 1365 -668 1399
rect -578 1365 -490 1399
rect -400 1365 -312 1399
rect -222 1365 -134 1399
rect -44 1365 44 1399
rect 134 1365 222 1399
rect 312 1365 400 1399
rect 490 1365 578 1399
rect 668 1365 756 1399
rect 846 1365 934 1399
rect 1024 1365 1112 1399
rect 1202 1365 1290 1399
rect 1380 1365 1468 1399
rect 1558 1365 1646 1399
rect 1736 1365 1824 1399
rect 1914 1365 2002 1399
rect 2092 1365 2180 1399
rect 2270 1365 2358 1399
rect 2448 1365 2536 1399
rect 2626 1365 2714 1399
rect 2804 1365 2892 1399
rect 2982 1365 3070 1399
rect 3160 1365 3248 1399
rect 3338 1365 3426 1399
rect 3516 1365 3604 1399
rect 3694 1365 3782 1399
rect 3872 1365 3960 1399
rect -4022 130 -3988 1306
rect -3844 130 -3810 1306
rect -3666 130 -3632 1306
rect -3488 130 -3454 1306
rect -3310 130 -3276 1306
rect -3132 130 -3098 1306
rect -2954 130 -2920 1306
rect -2776 130 -2742 1306
rect -2598 130 -2564 1306
rect -2420 130 -2386 1306
rect -2242 130 -2208 1306
rect -2064 130 -2030 1306
rect -1886 130 -1852 1306
rect -1708 130 -1674 1306
rect -1530 130 -1496 1306
rect -1352 130 -1318 1306
rect -1174 130 -1140 1306
rect -996 130 -962 1306
rect -818 130 -784 1306
rect -640 130 -606 1306
rect -462 130 -428 1306
rect -284 130 -250 1306
rect -106 130 -72 1306
rect 72 130 106 1306
rect 250 130 284 1306
rect 428 130 462 1306
rect 606 130 640 1306
rect 784 130 818 1306
rect 962 130 996 1306
rect 1140 130 1174 1306
rect 1318 130 1352 1306
rect 1496 130 1530 1306
rect 1674 130 1708 1306
rect 1852 130 1886 1306
rect 2030 130 2064 1306
rect 2208 130 2242 1306
rect 2386 130 2420 1306
rect 2564 130 2598 1306
rect 2742 130 2776 1306
rect 2920 130 2954 1306
rect 3098 130 3132 1306
rect 3276 130 3310 1306
rect 3454 130 3488 1306
rect 3632 130 3666 1306
rect 3810 130 3844 1306
rect 3988 130 4022 1306
rect -3960 37 -3872 71
rect -3782 37 -3694 71
rect -3604 37 -3516 71
rect -3426 37 -3338 71
rect -3248 37 -3160 71
rect -3070 37 -2982 71
rect -2892 37 -2804 71
rect -2714 37 -2626 71
rect -2536 37 -2448 71
rect -2358 37 -2270 71
rect -2180 37 -2092 71
rect -2002 37 -1914 71
rect -1824 37 -1736 71
rect -1646 37 -1558 71
rect -1468 37 -1380 71
rect -1290 37 -1202 71
rect -1112 37 -1024 71
rect -934 37 -846 71
rect -756 37 -668 71
rect -578 37 -490 71
rect -400 37 -312 71
rect -222 37 -134 71
rect -44 37 44 71
rect 134 37 222 71
rect 312 37 400 71
rect 490 37 578 71
rect 668 37 756 71
rect 846 37 934 71
rect 1024 37 1112 71
rect 1202 37 1290 71
rect 1380 37 1468 71
rect 1558 37 1646 71
rect 1736 37 1824 71
rect 1914 37 2002 71
rect 2092 37 2180 71
rect 2270 37 2358 71
rect 2448 37 2536 71
rect 2626 37 2714 71
rect 2804 37 2892 71
rect 2982 37 3070 71
rect 3160 37 3248 71
rect 3338 37 3426 71
rect 3516 37 3604 71
rect 3694 37 3782 71
rect 3872 37 3960 71
rect -3960 -71 -3872 -37
rect -3782 -71 -3694 -37
rect -3604 -71 -3516 -37
rect -3426 -71 -3338 -37
rect -3248 -71 -3160 -37
rect -3070 -71 -2982 -37
rect -2892 -71 -2804 -37
rect -2714 -71 -2626 -37
rect -2536 -71 -2448 -37
rect -2358 -71 -2270 -37
rect -2180 -71 -2092 -37
rect -2002 -71 -1914 -37
rect -1824 -71 -1736 -37
rect -1646 -71 -1558 -37
rect -1468 -71 -1380 -37
rect -1290 -71 -1202 -37
rect -1112 -71 -1024 -37
rect -934 -71 -846 -37
rect -756 -71 -668 -37
rect -578 -71 -490 -37
rect -400 -71 -312 -37
rect -222 -71 -134 -37
rect -44 -71 44 -37
rect 134 -71 222 -37
rect 312 -71 400 -37
rect 490 -71 578 -37
rect 668 -71 756 -37
rect 846 -71 934 -37
rect 1024 -71 1112 -37
rect 1202 -71 1290 -37
rect 1380 -71 1468 -37
rect 1558 -71 1646 -37
rect 1736 -71 1824 -37
rect 1914 -71 2002 -37
rect 2092 -71 2180 -37
rect 2270 -71 2358 -37
rect 2448 -71 2536 -37
rect 2626 -71 2714 -37
rect 2804 -71 2892 -37
rect 2982 -71 3070 -37
rect 3160 -71 3248 -37
rect 3338 -71 3426 -37
rect 3516 -71 3604 -37
rect 3694 -71 3782 -37
rect 3872 -71 3960 -37
rect -4022 -1306 -3988 -130
rect -3844 -1306 -3810 -130
rect -3666 -1306 -3632 -130
rect -3488 -1306 -3454 -130
rect -3310 -1306 -3276 -130
rect -3132 -1306 -3098 -130
rect -2954 -1306 -2920 -130
rect -2776 -1306 -2742 -130
rect -2598 -1306 -2564 -130
rect -2420 -1306 -2386 -130
rect -2242 -1306 -2208 -130
rect -2064 -1306 -2030 -130
rect -1886 -1306 -1852 -130
rect -1708 -1306 -1674 -130
rect -1530 -1306 -1496 -130
rect -1352 -1306 -1318 -130
rect -1174 -1306 -1140 -130
rect -996 -1306 -962 -130
rect -818 -1306 -784 -130
rect -640 -1306 -606 -130
rect -462 -1306 -428 -130
rect -284 -1306 -250 -130
rect -106 -1306 -72 -130
rect 72 -1306 106 -130
rect 250 -1306 284 -130
rect 428 -1306 462 -130
rect 606 -1306 640 -130
rect 784 -1306 818 -130
rect 962 -1306 996 -130
rect 1140 -1306 1174 -130
rect 1318 -1306 1352 -130
rect 1496 -1306 1530 -130
rect 1674 -1306 1708 -130
rect 1852 -1306 1886 -130
rect 2030 -1306 2064 -130
rect 2208 -1306 2242 -130
rect 2386 -1306 2420 -130
rect 2564 -1306 2598 -130
rect 2742 -1306 2776 -130
rect 2920 -1306 2954 -130
rect 3098 -1306 3132 -130
rect 3276 -1306 3310 -130
rect 3454 -1306 3488 -130
rect 3632 -1306 3666 -130
rect 3810 -1306 3844 -130
rect 3988 -1306 4022 -130
rect -3960 -1399 -3872 -1365
rect -3782 -1399 -3694 -1365
rect -3604 -1399 -3516 -1365
rect -3426 -1399 -3338 -1365
rect -3248 -1399 -3160 -1365
rect -3070 -1399 -2982 -1365
rect -2892 -1399 -2804 -1365
rect -2714 -1399 -2626 -1365
rect -2536 -1399 -2448 -1365
rect -2358 -1399 -2270 -1365
rect -2180 -1399 -2092 -1365
rect -2002 -1399 -1914 -1365
rect -1824 -1399 -1736 -1365
rect -1646 -1399 -1558 -1365
rect -1468 -1399 -1380 -1365
rect -1290 -1399 -1202 -1365
rect -1112 -1399 -1024 -1365
rect -934 -1399 -846 -1365
rect -756 -1399 -668 -1365
rect -578 -1399 -490 -1365
rect -400 -1399 -312 -1365
rect -222 -1399 -134 -1365
rect -44 -1399 44 -1365
rect 134 -1399 222 -1365
rect 312 -1399 400 -1365
rect 490 -1399 578 -1365
rect 668 -1399 756 -1365
rect 846 -1399 934 -1365
rect 1024 -1399 1112 -1365
rect 1202 -1399 1290 -1365
rect 1380 -1399 1468 -1365
rect 1558 -1399 1646 -1365
rect 1736 -1399 1824 -1365
rect 1914 -1399 2002 -1365
rect 2092 -1399 2180 -1365
rect 2270 -1399 2358 -1365
rect 2448 -1399 2536 -1365
rect 2626 -1399 2714 -1365
rect 2804 -1399 2892 -1365
rect 2982 -1399 3070 -1365
rect 3160 -1399 3248 -1365
rect 3338 -1399 3426 -1365
rect 3516 -1399 3604 -1365
rect 3694 -1399 3782 -1365
rect 3872 -1399 3960 -1365
<< metal1 >>
rect -3972 1399 -3860 1405
rect -3972 1365 -3960 1399
rect -3872 1365 -3860 1399
rect -3972 1359 -3860 1365
rect -3794 1399 -3682 1405
rect -3794 1365 -3782 1399
rect -3694 1365 -3682 1399
rect -3794 1359 -3682 1365
rect -3616 1399 -3504 1405
rect -3616 1365 -3604 1399
rect -3516 1365 -3504 1399
rect -3616 1359 -3504 1365
rect -3438 1399 -3326 1405
rect -3438 1365 -3426 1399
rect -3338 1365 -3326 1399
rect -3438 1359 -3326 1365
rect -3260 1399 -3148 1405
rect -3260 1365 -3248 1399
rect -3160 1365 -3148 1399
rect -3260 1359 -3148 1365
rect -3082 1399 -2970 1405
rect -3082 1365 -3070 1399
rect -2982 1365 -2970 1399
rect -3082 1359 -2970 1365
rect -2904 1399 -2792 1405
rect -2904 1365 -2892 1399
rect -2804 1365 -2792 1399
rect -2904 1359 -2792 1365
rect -2726 1399 -2614 1405
rect -2726 1365 -2714 1399
rect -2626 1365 -2614 1399
rect -2726 1359 -2614 1365
rect -2548 1399 -2436 1405
rect -2548 1365 -2536 1399
rect -2448 1365 -2436 1399
rect -2548 1359 -2436 1365
rect -2370 1399 -2258 1405
rect -2370 1365 -2358 1399
rect -2270 1365 -2258 1399
rect -2370 1359 -2258 1365
rect -2192 1399 -2080 1405
rect -2192 1365 -2180 1399
rect -2092 1365 -2080 1399
rect -2192 1359 -2080 1365
rect -2014 1399 -1902 1405
rect -2014 1365 -2002 1399
rect -1914 1365 -1902 1399
rect -2014 1359 -1902 1365
rect -1836 1399 -1724 1405
rect -1836 1365 -1824 1399
rect -1736 1365 -1724 1399
rect -1836 1359 -1724 1365
rect -1658 1399 -1546 1405
rect -1658 1365 -1646 1399
rect -1558 1365 -1546 1399
rect -1658 1359 -1546 1365
rect -1480 1399 -1368 1405
rect -1480 1365 -1468 1399
rect -1380 1365 -1368 1399
rect -1480 1359 -1368 1365
rect -1302 1399 -1190 1405
rect -1302 1365 -1290 1399
rect -1202 1365 -1190 1399
rect -1302 1359 -1190 1365
rect -1124 1399 -1012 1405
rect -1124 1365 -1112 1399
rect -1024 1365 -1012 1399
rect -1124 1359 -1012 1365
rect -946 1399 -834 1405
rect -946 1365 -934 1399
rect -846 1365 -834 1399
rect -946 1359 -834 1365
rect -768 1399 -656 1405
rect -768 1365 -756 1399
rect -668 1365 -656 1399
rect -768 1359 -656 1365
rect -590 1399 -478 1405
rect -590 1365 -578 1399
rect -490 1365 -478 1399
rect -590 1359 -478 1365
rect -412 1399 -300 1405
rect -412 1365 -400 1399
rect -312 1365 -300 1399
rect -412 1359 -300 1365
rect -234 1399 -122 1405
rect -234 1365 -222 1399
rect -134 1365 -122 1399
rect -234 1359 -122 1365
rect -56 1399 56 1405
rect -56 1365 -44 1399
rect 44 1365 56 1399
rect -56 1359 56 1365
rect 122 1399 234 1405
rect 122 1365 134 1399
rect 222 1365 234 1399
rect 122 1359 234 1365
rect 300 1399 412 1405
rect 300 1365 312 1399
rect 400 1365 412 1399
rect 300 1359 412 1365
rect 478 1399 590 1405
rect 478 1365 490 1399
rect 578 1365 590 1399
rect 478 1359 590 1365
rect 656 1399 768 1405
rect 656 1365 668 1399
rect 756 1365 768 1399
rect 656 1359 768 1365
rect 834 1399 946 1405
rect 834 1365 846 1399
rect 934 1365 946 1399
rect 834 1359 946 1365
rect 1012 1399 1124 1405
rect 1012 1365 1024 1399
rect 1112 1365 1124 1399
rect 1012 1359 1124 1365
rect 1190 1399 1302 1405
rect 1190 1365 1202 1399
rect 1290 1365 1302 1399
rect 1190 1359 1302 1365
rect 1368 1399 1480 1405
rect 1368 1365 1380 1399
rect 1468 1365 1480 1399
rect 1368 1359 1480 1365
rect 1546 1399 1658 1405
rect 1546 1365 1558 1399
rect 1646 1365 1658 1399
rect 1546 1359 1658 1365
rect 1724 1399 1836 1405
rect 1724 1365 1736 1399
rect 1824 1365 1836 1399
rect 1724 1359 1836 1365
rect 1902 1399 2014 1405
rect 1902 1365 1914 1399
rect 2002 1365 2014 1399
rect 1902 1359 2014 1365
rect 2080 1399 2192 1405
rect 2080 1365 2092 1399
rect 2180 1365 2192 1399
rect 2080 1359 2192 1365
rect 2258 1399 2370 1405
rect 2258 1365 2270 1399
rect 2358 1365 2370 1399
rect 2258 1359 2370 1365
rect 2436 1399 2548 1405
rect 2436 1365 2448 1399
rect 2536 1365 2548 1399
rect 2436 1359 2548 1365
rect 2614 1399 2726 1405
rect 2614 1365 2626 1399
rect 2714 1365 2726 1399
rect 2614 1359 2726 1365
rect 2792 1399 2904 1405
rect 2792 1365 2804 1399
rect 2892 1365 2904 1399
rect 2792 1359 2904 1365
rect 2970 1399 3082 1405
rect 2970 1365 2982 1399
rect 3070 1365 3082 1399
rect 2970 1359 3082 1365
rect 3148 1399 3260 1405
rect 3148 1365 3160 1399
rect 3248 1365 3260 1399
rect 3148 1359 3260 1365
rect 3326 1399 3438 1405
rect 3326 1365 3338 1399
rect 3426 1365 3438 1399
rect 3326 1359 3438 1365
rect 3504 1399 3616 1405
rect 3504 1365 3516 1399
rect 3604 1365 3616 1399
rect 3504 1359 3616 1365
rect 3682 1399 3794 1405
rect 3682 1365 3694 1399
rect 3782 1365 3794 1399
rect 3682 1359 3794 1365
rect 3860 1399 3972 1405
rect 3860 1365 3872 1399
rect 3960 1365 3972 1399
rect 3860 1359 3972 1365
rect -4028 1306 -3982 1318
rect -4028 130 -4022 1306
rect -3988 130 -3982 1306
rect -4028 118 -3982 130
rect -3850 1306 -3804 1318
rect -3850 130 -3844 1306
rect -3810 130 -3804 1306
rect -3850 118 -3804 130
rect -3672 1306 -3626 1318
rect -3672 130 -3666 1306
rect -3632 130 -3626 1306
rect -3672 118 -3626 130
rect -3494 1306 -3448 1318
rect -3494 130 -3488 1306
rect -3454 130 -3448 1306
rect -3494 118 -3448 130
rect -3316 1306 -3270 1318
rect -3316 130 -3310 1306
rect -3276 130 -3270 1306
rect -3316 118 -3270 130
rect -3138 1306 -3092 1318
rect -3138 130 -3132 1306
rect -3098 130 -3092 1306
rect -3138 118 -3092 130
rect -2960 1306 -2914 1318
rect -2960 130 -2954 1306
rect -2920 130 -2914 1306
rect -2960 118 -2914 130
rect -2782 1306 -2736 1318
rect -2782 130 -2776 1306
rect -2742 130 -2736 1306
rect -2782 118 -2736 130
rect -2604 1306 -2558 1318
rect -2604 130 -2598 1306
rect -2564 130 -2558 1306
rect -2604 118 -2558 130
rect -2426 1306 -2380 1318
rect -2426 130 -2420 1306
rect -2386 130 -2380 1306
rect -2426 118 -2380 130
rect -2248 1306 -2202 1318
rect -2248 130 -2242 1306
rect -2208 130 -2202 1306
rect -2248 118 -2202 130
rect -2070 1306 -2024 1318
rect -2070 130 -2064 1306
rect -2030 130 -2024 1306
rect -2070 118 -2024 130
rect -1892 1306 -1846 1318
rect -1892 130 -1886 1306
rect -1852 130 -1846 1306
rect -1892 118 -1846 130
rect -1714 1306 -1668 1318
rect -1714 130 -1708 1306
rect -1674 130 -1668 1306
rect -1714 118 -1668 130
rect -1536 1306 -1490 1318
rect -1536 130 -1530 1306
rect -1496 130 -1490 1306
rect -1536 118 -1490 130
rect -1358 1306 -1312 1318
rect -1358 130 -1352 1306
rect -1318 130 -1312 1306
rect -1358 118 -1312 130
rect -1180 1306 -1134 1318
rect -1180 130 -1174 1306
rect -1140 130 -1134 1306
rect -1180 118 -1134 130
rect -1002 1306 -956 1318
rect -1002 130 -996 1306
rect -962 130 -956 1306
rect -1002 118 -956 130
rect -824 1306 -778 1318
rect -824 130 -818 1306
rect -784 130 -778 1306
rect -824 118 -778 130
rect -646 1306 -600 1318
rect -646 130 -640 1306
rect -606 130 -600 1306
rect -646 118 -600 130
rect -468 1306 -422 1318
rect -468 130 -462 1306
rect -428 130 -422 1306
rect -468 118 -422 130
rect -290 1306 -244 1318
rect -290 130 -284 1306
rect -250 130 -244 1306
rect -290 118 -244 130
rect -112 1306 -66 1318
rect -112 130 -106 1306
rect -72 130 -66 1306
rect -112 118 -66 130
rect 66 1306 112 1318
rect 66 130 72 1306
rect 106 130 112 1306
rect 66 118 112 130
rect 244 1306 290 1318
rect 244 130 250 1306
rect 284 130 290 1306
rect 244 118 290 130
rect 422 1306 468 1318
rect 422 130 428 1306
rect 462 130 468 1306
rect 422 118 468 130
rect 600 1306 646 1318
rect 600 130 606 1306
rect 640 130 646 1306
rect 600 118 646 130
rect 778 1306 824 1318
rect 778 130 784 1306
rect 818 130 824 1306
rect 778 118 824 130
rect 956 1306 1002 1318
rect 956 130 962 1306
rect 996 130 1002 1306
rect 956 118 1002 130
rect 1134 1306 1180 1318
rect 1134 130 1140 1306
rect 1174 130 1180 1306
rect 1134 118 1180 130
rect 1312 1306 1358 1318
rect 1312 130 1318 1306
rect 1352 130 1358 1306
rect 1312 118 1358 130
rect 1490 1306 1536 1318
rect 1490 130 1496 1306
rect 1530 130 1536 1306
rect 1490 118 1536 130
rect 1668 1306 1714 1318
rect 1668 130 1674 1306
rect 1708 130 1714 1306
rect 1668 118 1714 130
rect 1846 1306 1892 1318
rect 1846 130 1852 1306
rect 1886 130 1892 1306
rect 1846 118 1892 130
rect 2024 1306 2070 1318
rect 2024 130 2030 1306
rect 2064 130 2070 1306
rect 2024 118 2070 130
rect 2202 1306 2248 1318
rect 2202 130 2208 1306
rect 2242 130 2248 1306
rect 2202 118 2248 130
rect 2380 1306 2426 1318
rect 2380 130 2386 1306
rect 2420 130 2426 1306
rect 2380 118 2426 130
rect 2558 1306 2604 1318
rect 2558 130 2564 1306
rect 2598 130 2604 1306
rect 2558 118 2604 130
rect 2736 1306 2782 1318
rect 2736 130 2742 1306
rect 2776 130 2782 1306
rect 2736 118 2782 130
rect 2914 1306 2960 1318
rect 2914 130 2920 1306
rect 2954 130 2960 1306
rect 2914 118 2960 130
rect 3092 1306 3138 1318
rect 3092 130 3098 1306
rect 3132 130 3138 1306
rect 3092 118 3138 130
rect 3270 1306 3316 1318
rect 3270 130 3276 1306
rect 3310 130 3316 1306
rect 3270 118 3316 130
rect 3448 1306 3494 1318
rect 3448 130 3454 1306
rect 3488 130 3494 1306
rect 3448 118 3494 130
rect 3626 1306 3672 1318
rect 3626 130 3632 1306
rect 3666 130 3672 1306
rect 3626 118 3672 130
rect 3804 1306 3850 1318
rect 3804 130 3810 1306
rect 3844 130 3850 1306
rect 3804 118 3850 130
rect 3982 1306 4028 1318
rect 3982 130 3988 1306
rect 4022 130 4028 1306
rect 3982 118 4028 130
rect -3972 71 -3860 77
rect -3972 37 -3960 71
rect -3872 37 -3860 71
rect -3972 31 -3860 37
rect -3794 71 -3682 77
rect -3794 37 -3782 71
rect -3694 37 -3682 71
rect -3794 31 -3682 37
rect -3616 71 -3504 77
rect -3616 37 -3604 71
rect -3516 37 -3504 71
rect -3616 31 -3504 37
rect -3438 71 -3326 77
rect -3438 37 -3426 71
rect -3338 37 -3326 71
rect -3438 31 -3326 37
rect -3260 71 -3148 77
rect -3260 37 -3248 71
rect -3160 37 -3148 71
rect -3260 31 -3148 37
rect -3082 71 -2970 77
rect -3082 37 -3070 71
rect -2982 37 -2970 71
rect -3082 31 -2970 37
rect -2904 71 -2792 77
rect -2904 37 -2892 71
rect -2804 37 -2792 71
rect -2904 31 -2792 37
rect -2726 71 -2614 77
rect -2726 37 -2714 71
rect -2626 37 -2614 71
rect -2726 31 -2614 37
rect -2548 71 -2436 77
rect -2548 37 -2536 71
rect -2448 37 -2436 71
rect -2548 31 -2436 37
rect -2370 71 -2258 77
rect -2370 37 -2358 71
rect -2270 37 -2258 71
rect -2370 31 -2258 37
rect -2192 71 -2080 77
rect -2192 37 -2180 71
rect -2092 37 -2080 71
rect -2192 31 -2080 37
rect -2014 71 -1902 77
rect -2014 37 -2002 71
rect -1914 37 -1902 71
rect -2014 31 -1902 37
rect -1836 71 -1724 77
rect -1836 37 -1824 71
rect -1736 37 -1724 71
rect -1836 31 -1724 37
rect -1658 71 -1546 77
rect -1658 37 -1646 71
rect -1558 37 -1546 71
rect -1658 31 -1546 37
rect -1480 71 -1368 77
rect -1480 37 -1468 71
rect -1380 37 -1368 71
rect -1480 31 -1368 37
rect -1302 71 -1190 77
rect -1302 37 -1290 71
rect -1202 37 -1190 71
rect -1302 31 -1190 37
rect -1124 71 -1012 77
rect -1124 37 -1112 71
rect -1024 37 -1012 71
rect -1124 31 -1012 37
rect -946 71 -834 77
rect -946 37 -934 71
rect -846 37 -834 71
rect -946 31 -834 37
rect -768 71 -656 77
rect -768 37 -756 71
rect -668 37 -656 71
rect -768 31 -656 37
rect -590 71 -478 77
rect -590 37 -578 71
rect -490 37 -478 71
rect -590 31 -478 37
rect -412 71 -300 77
rect -412 37 -400 71
rect -312 37 -300 71
rect -412 31 -300 37
rect -234 71 -122 77
rect -234 37 -222 71
rect -134 37 -122 71
rect -234 31 -122 37
rect -56 71 56 77
rect -56 37 -44 71
rect 44 37 56 71
rect -56 31 56 37
rect 122 71 234 77
rect 122 37 134 71
rect 222 37 234 71
rect 122 31 234 37
rect 300 71 412 77
rect 300 37 312 71
rect 400 37 412 71
rect 300 31 412 37
rect 478 71 590 77
rect 478 37 490 71
rect 578 37 590 71
rect 478 31 590 37
rect 656 71 768 77
rect 656 37 668 71
rect 756 37 768 71
rect 656 31 768 37
rect 834 71 946 77
rect 834 37 846 71
rect 934 37 946 71
rect 834 31 946 37
rect 1012 71 1124 77
rect 1012 37 1024 71
rect 1112 37 1124 71
rect 1012 31 1124 37
rect 1190 71 1302 77
rect 1190 37 1202 71
rect 1290 37 1302 71
rect 1190 31 1302 37
rect 1368 71 1480 77
rect 1368 37 1380 71
rect 1468 37 1480 71
rect 1368 31 1480 37
rect 1546 71 1658 77
rect 1546 37 1558 71
rect 1646 37 1658 71
rect 1546 31 1658 37
rect 1724 71 1836 77
rect 1724 37 1736 71
rect 1824 37 1836 71
rect 1724 31 1836 37
rect 1902 71 2014 77
rect 1902 37 1914 71
rect 2002 37 2014 71
rect 1902 31 2014 37
rect 2080 71 2192 77
rect 2080 37 2092 71
rect 2180 37 2192 71
rect 2080 31 2192 37
rect 2258 71 2370 77
rect 2258 37 2270 71
rect 2358 37 2370 71
rect 2258 31 2370 37
rect 2436 71 2548 77
rect 2436 37 2448 71
rect 2536 37 2548 71
rect 2436 31 2548 37
rect 2614 71 2726 77
rect 2614 37 2626 71
rect 2714 37 2726 71
rect 2614 31 2726 37
rect 2792 71 2904 77
rect 2792 37 2804 71
rect 2892 37 2904 71
rect 2792 31 2904 37
rect 2970 71 3082 77
rect 2970 37 2982 71
rect 3070 37 3082 71
rect 2970 31 3082 37
rect 3148 71 3260 77
rect 3148 37 3160 71
rect 3248 37 3260 71
rect 3148 31 3260 37
rect 3326 71 3438 77
rect 3326 37 3338 71
rect 3426 37 3438 71
rect 3326 31 3438 37
rect 3504 71 3616 77
rect 3504 37 3516 71
rect 3604 37 3616 71
rect 3504 31 3616 37
rect 3682 71 3794 77
rect 3682 37 3694 71
rect 3782 37 3794 71
rect 3682 31 3794 37
rect 3860 71 3972 77
rect 3860 37 3872 71
rect 3960 37 3972 71
rect 3860 31 3972 37
rect -3972 -37 -3860 -31
rect -3972 -71 -3960 -37
rect -3872 -71 -3860 -37
rect -3972 -77 -3860 -71
rect -3794 -37 -3682 -31
rect -3794 -71 -3782 -37
rect -3694 -71 -3682 -37
rect -3794 -77 -3682 -71
rect -3616 -37 -3504 -31
rect -3616 -71 -3604 -37
rect -3516 -71 -3504 -37
rect -3616 -77 -3504 -71
rect -3438 -37 -3326 -31
rect -3438 -71 -3426 -37
rect -3338 -71 -3326 -37
rect -3438 -77 -3326 -71
rect -3260 -37 -3148 -31
rect -3260 -71 -3248 -37
rect -3160 -71 -3148 -37
rect -3260 -77 -3148 -71
rect -3082 -37 -2970 -31
rect -3082 -71 -3070 -37
rect -2982 -71 -2970 -37
rect -3082 -77 -2970 -71
rect -2904 -37 -2792 -31
rect -2904 -71 -2892 -37
rect -2804 -71 -2792 -37
rect -2904 -77 -2792 -71
rect -2726 -37 -2614 -31
rect -2726 -71 -2714 -37
rect -2626 -71 -2614 -37
rect -2726 -77 -2614 -71
rect -2548 -37 -2436 -31
rect -2548 -71 -2536 -37
rect -2448 -71 -2436 -37
rect -2548 -77 -2436 -71
rect -2370 -37 -2258 -31
rect -2370 -71 -2358 -37
rect -2270 -71 -2258 -37
rect -2370 -77 -2258 -71
rect -2192 -37 -2080 -31
rect -2192 -71 -2180 -37
rect -2092 -71 -2080 -37
rect -2192 -77 -2080 -71
rect -2014 -37 -1902 -31
rect -2014 -71 -2002 -37
rect -1914 -71 -1902 -37
rect -2014 -77 -1902 -71
rect -1836 -37 -1724 -31
rect -1836 -71 -1824 -37
rect -1736 -71 -1724 -37
rect -1836 -77 -1724 -71
rect -1658 -37 -1546 -31
rect -1658 -71 -1646 -37
rect -1558 -71 -1546 -37
rect -1658 -77 -1546 -71
rect -1480 -37 -1368 -31
rect -1480 -71 -1468 -37
rect -1380 -71 -1368 -37
rect -1480 -77 -1368 -71
rect -1302 -37 -1190 -31
rect -1302 -71 -1290 -37
rect -1202 -71 -1190 -37
rect -1302 -77 -1190 -71
rect -1124 -37 -1012 -31
rect -1124 -71 -1112 -37
rect -1024 -71 -1012 -37
rect -1124 -77 -1012 -71
rect -946 -37 -834 -31
rect -946 -71 -934 -37
rect -846 -71 -834 -37
rect -946 -77 -834 -71
rect -768 -37 -656 -31
rect -768 -71 -756 -37
rect -668 -71 -656 -37
rect -768 -77 -656 -71
rect -590 -37 -478 -31
rect -590 -71 -578 -37
rect -490 -71 -478 -37
rect -590 -77 -478 -71
rect -412 -37 -300 -31
rect -412 -71 -400 -37
rect -312 -71 -300 -37
rect -412 -77 -300 -71
rect -234 -37 -122 -31
rect -234 -71 -222 -37
rect -134 -71 -122 -37
rect -234 -77 -122 -71
rect -56 -37 56 -31
rect -56 -71 -44 -37
rect 44 -71 56 -37
rect -56 -77 56 -71
rect 122 -37 234 -31
rect 122 -71 134 -37
rect 222 -71 234 -37
rect 122 -77 234 -71
rect 300 -37 412 -31
rect 300 -71 312 -37
rect 400 -71 412 -37
rect 300 -77 412 -71
rect 478 -37 590 -31
rect 478 -71 490 -37
rect 578 -71 590 -37
rect 478 -77 590 -71
rect 656 -37 768 -31
rect 656 -71 668 -37
rect 756 -71 768 -37
rect 656 -77 768 -71
rect 834 -37 946 -31
rect 834 -71 846 -37
rect 934 -71 946 -37
rect 834 -77 946 -71
rect 1012 -37 1124 -31
rect 1012 -71 1024 -37
rect 1112 -71 1124 -37
rect 1012 -77 1124 -71
rect 1190 -37 1302 -31
rect 1190 -71 1202 -37
rect 1290 -71 1302 -37
rect 1190 -77 1302 -71
rect 1368 -37 1480 -31
rect 1368 -71 1380 -37
rect 1468 -71 1480 -37
rect 1368 -77 1480 -71
rect 1546 -37 1658 -31
rect 1546 -71 1558 -37
rect 1646 -71 1658 -37
rect 1546 -77 1658 -71
rect 1724 -37 1836 -31
rect 1724 -71 1736 -37
rect 1824 -71 1836 -37
rect 1724 -77 1836 -71
rect 1902 -37 2014 -31
rect 1902 -71 1914 -37
rect 2002 -71 2014 -37
rect 1902 -77 2014 -71
rect 2080 -37 2192 -31
rect 2080 -71 2092 -37
rect 2180 -71 2192 -37
rect 2080 -77 2192 -71
rect 2258 -37 2370 -31
rect 2258 -71 2270 -37
rect 2358 -71 2370 -37
rect 2258 -77 2370 -71
rect 2436 -37 2548 -31
rect 2436 -71 2448 -37
rect 2536 -71 2548 -37
rect 2436 -77 2548 -71
rect 2614 -37 2726 -31
rect 2614 -71 2626 -37
rect 2714 -71 2726 -37
rect 2614 -77 2726 -71
rect 2792 -37 2904 -31
rect 2792 -71 2804 -37
rect 2892 -71 2904 -37
rect 2792 -77 2904 -71
rect 2970 -37 3082 -31
rect 2970 -71 2982 -37
rect 3070 -71 3082 -37
rect 2970 -77 3082 -71
rect 3148 -37 3260 -31
rect 3148 -71 3160 -37
rect 3248 -71 3260 -37
rect 3148 -77 3260 -71
rect 3326 -37 3438 -31
rect 3326 -71 3338 -37
rect 3426 -71 3438 -37
rect 3326 -77 3438 -71
rect 3504 -37 3616 -31
rect 3504 -71 3516 -37
rect 3604 -71 3616 -37
rect 3504 -77 3616 -71
rect 3682 -37 3794 -31
rect 3682 -71 3694 -37
rect 3782 -71 3794 -37
rect 3682 -77 3794 -71
rect 3860 -37 3972 -31
rect 3860 -71 3872 -37
rect 3960 -71 3972 -37
rect 3860 -77 3972 -71
rect -4028 -130 -3982 -118
rect -4028 -1306 -4022 -130
rect -3988 -1306 -3982 -130
rect -4028 -1318 -3982 -1306
rect -3850 -130 -3804 -118
rect -3850 -1306 -3844 -130
rect -3810 -1306 -3804 -130
rect -3850 -1318 -3804 -1306
rect -3672 -130 -3626 -118
rect -3672 -1306 -3666 -130
rect -3632 -1306 -3626 -130
rect -3672 -1318 -3626 -1306
rect -3494 -130 -3448 -118
rect -3494 -1306 -3488 -130
rect -3454 -1306 -3448 -130
rect -3494 -1318 -3448 -1306
rect -3316 -130 -3270 -118
rect -3316 -1306 -3310 -130
rect -3276 -1306 -3270 -130
rect -3316 -1318 -3270 -1306
rect -3138 -130 -3092 -118
rect -3138 -1306 -3132 -130
rect -3098 -1306 -3092 -130
rect -3138 -1318 -3092 -1306
rect -2960 -130 -2914 -118
rect -2960 -1306 -2954 -130
rect -2920 -1306 -2914 -130
rect -2960 -1318 -2914 -1306
rect -2782 -130 -2736 -118
rect -2782 -1306 -2776 -130
rect -2742 -1306 -2736 -130
rect -2782 -1318 -2736 -1306
rect -2604 -130 -2558 -118
rect -2604 -1306 -2598 -130
rect -2564 -1306 -2558 -130
rect -2604 -1318 -2558 -1306
rect -2426 -130 -2380 -118
rect -2426 -1306 -2420 -130
rect -2386 -1306 -2380 -130
rect -2426 -1318 -2380 -1306
rect -2248 -130 -2202 -118
rect -2248 -1306 -2242 -130
rect -2208 -1306 -2202 -130
rect -2248 -1318 -2202 -1306
rect -2070 -130 -2024 -118
rect -2070 -1306 -2064 -130
rect -2030 -1306 -2024 -130
rect -2070 -1318 -2024 -1306
rect -1892 -130 -1846 -118
rect -1892 -1306 -1886 -130
rect -1852 -1306 -1846 -130
rect -1892 -1318 -1846 -1306
rect -1714 -130 -1668 -118
rect -1714 -1306 -1708 -130
rect -1674 -1306 -1668 -130
rect -1714 -1318 -1668 -1306
rect -1536 -130 -1490 -118
rect -1536 -1306 -1530 -130
rect -1496 -1306 -1490 -130
rect -1536 -1318 -1490 -1306
rect -1358 -130 -1312 -118
rect -1358 -1306 -1352 -130
rect -1318 -1306 -1312 -130
rect -1358 -1318 -1312 -1306
rect -1180 -130 -1134 -118
rect -1180 -1306 -1174 -130
rect -1140 -1306 -1134 -130
rect -1180 -1318 -1134 -1306
rect -1002 -130 -956 -118
rect -1002 -1306 -996 -130
rect -962 -1306 -956 -130
rect -1002 -1318 -956 -1306
rect -824 -130 -778 -118
rect -824 -1306 -818 -130
rect -784 -1306 -778 -130
rect -824 -1318 -778 -1306
rect -646 -130 -600 -118
rect -646 -1306 -640 -130
rect -606 -1306 -600 -130
rect -646 -1318 -600 -1306
rect -468 -130 -422 -118
rect -468 -1306 -462 -130
rect -428 -1306 -422 -130
rect -468 -1318 -422 -1306
rect -290 -130 -244 -118
rect -290 -1306 -284 -130
rect -250 -1306 -244 -130
rect -290 -1318 -244 -1306
rect -112 -130 -66 -118
rect -112 -1306 -106 -130
rect -72 -1306 -66 -130
rect -112 -1318 -66 -1306
rect 66 -130 112 -118
rect 66 -1306 72 -130
rect 106 -1306 112 -130
rect 66 -1318 112 -1306
rect 244 -130 290 -118
rect 244 -1306 250 -130
rect 284 -1306 290 -130
rect 244 -1318 290 -1306
rect 422 -130 468 -118
rect 422 -1306 428 -130
rect 462 -1306 468 -130
rect 422 -1318 468 -1306
rect 600 -130 646 -118
rect 600 -1306 606 -130
rect 640 -1306 646 -130
rect 600 -1318 646 -1306
rect 778 -130 824 -118
rect 778 -1306 784 -130
rect 818 -1306 824 -130
rect 778 -1318 824 -1306
rect 956 -130 1002 -118
rect 956 -1306 962 -130
rect 996 -1306 1002 -130
rect 956 -1318 1002 -1306
rect 1134 -130 1180 -118
rect 1134 -1306 1140 -130
rect 1174 -1306 1180 -130
rect 1134 -1318 1180 -1306
rect 1312 -130 1358 -118
rect 1312 -1306 1318 -130
rect 1352 -1306 1358 -130
rect 1312 -1318 1358 -1306
rect 1490 -130 1536 -118
rect 1490 -1306 1496 -130
rect 1530 -1306 1536 -130
rect 1490 -1318 1536 -1306
rect 1668 -130 1714 -118
rect 1668 -1306 1674 -130
rect 1708 -1306 1714 -130
rect 1668 -1318 1714 -1306
rect 1846 -130 1892 -118
rect 1846 -1306 1852 -130
rect 1886 -1306 1892 -130
rect 1846 -1318 1892 -1306
rect 2024 -130 2070 -118
rect 2024 -1306 2030 -130
rect 2064 -1306 2070 -130
rect 2024 -1318 2070 -1306
rect 2202 -130 2248 -118
rect 2202 -1306 2208 -130
rect 2242 -1306 2248 -130
rect 2202 -1318 2248 -1306
rect 2380 -130 2426 -118
rect 2380 -1306 2386 -130
rect 2420 -1306 2426 -130
rect 2380 -1318 2426 -1306
rect 2558 -130 2604 -118
rect 2558 -1306 2564 -130
rect 2598 -1306 2604 -130
rect 2558 -1318 2604 -1306
rect 2736 -130 2782 -118
rect 2736 -1306 2742 -130
rect 2776 -1306 2782 -130
rect 2736 -1318 2782 -1306
rect 2914 -130 2960 -118
rect 2914 -1306 2920 -130
rect 2954 -1306 2960 -130
rect 2914 -1318 2960 -1306
rect 3092 -130 3138 -118
rect 3092 -1306 3098 -130
rect 3132 -1306 3138 -130
rect 3092 -1318 3138 -1306
rect 3270 -130 3316 -118
rect 3270 -1306 3276 -130
rect 3310 -1306 3316 -130
rect 3270 -1318 3316 -1306
rect 3448 -130 3494 -118
rect 3448 -1306 3454 -130
rect 3488 -1306 3494 -130
rect 3448 -1318 3494 -1306
rect 3626 -130 3672 -118
rect 3626 -1306 3632 -130
rect 3666 -1306 3672 -130
rect 3626 -1318 3672 -1306
rect 3804 -130 3850 -118
rect 3804 -1306 3810 -130
rect 3844 -1306 3850 -130
rect 3804 -1318 3850 -1306
rect 3982 -130 4028 -118
rect 3982 -1306 3988 -130
rect 4022 -1306 4028 -130
rect 3982 -1318 4028 -1306
rect -3972 -1365 -3860 -1359
rect -3972 -1399 -3960 -1365
rect -3872 -1399 -3860 -1365
rect -3972 -1405 -3860 -1399
rect -3794 -1365 -3682 -1359
rect -3794 -1399 -3782 -1365
rect -3694 -1399 -3682 -1365
rect -3794 -1405 -3682 -1399
rect -3616 -1365 -3504 -1359
rect -3616 -1399 -3604 -1365
rect -3516 -1399 -3504 -1365
rect -3616 -1405 -3504 -1399
rect -3438 -1365 -3326 -1359
rect -3438 -1399 -3426 -1365
rect -3338 -1399 -3326 -1365
rect -3438 -1405 -3326 -1399
rect -3260 -1365 -3148 -1359
rect -3260 -1399 -3248 -1365
rect -3160 -1399 -3148 -1365
rect -3260 -1405 -3148 -1399
rect -3082 -1365 -2970 -1359
rect -3082 -1399 -3070 -1365
rect -2982 -1399 -2970 -1365
rect -3082 -1405 -2970 -1399
rect -2904 -1365 -2792 -1359
rect -2904 -1399 -2892 -1365
rect -2804 -1399 -2792 -1365
rect -2904 -1405 -2792 -1399
rect -2726 -1365 -2614 -1359
rect -2726 -1399 -2714 -1365
rect -2626 -1399 -2614 -1365
rect -2726 -1405 -2614 -1399
rect -2548 -1365 -2436 -1359
rect -2548 -1399 -2536 -1365
rect -2448 -1399 -2436 -1365
rect -2548 -1405 -2436 -1399
rect -2370 -1365 -2258 -1359
rect -2370 -1399 -2358 -1365
rect -2270 -1399 -2258 -1365
rect -2370 -1405 -2258 -1399
rect -2192 -1365 -2080 -1359
rect -2192 -1399 -2180 -1365
rect -2092 -1399 -2080 -1365
rect -2192 -1405 -2080 -1399
rect -2014 -1365 -1902 -1359
rect -2014 -1399 -2002 -1365
rect -1914 -1399 -1902 -1365
rect -2014 -1405 -1902 -1399
rect -1836 -1365 -1724 -1359
rect -1836 -1399 -1824 -1365
rect -1736 -1399 -1724 -1365
rect -1836 -1405 -1724 -1399
rect -1658 -1365 -1546 -1359
rect -1658 -1399 -1646 -1365
rect -1558 -1399 -1546 -1365
rect -1658 -1405 -1546 -1399
rect -1480 -1365 -1368 -1359
rect -1480 -1399 -1468 -1365
rect -1380 -1399 -1368 -1365
rect -1480 -1405 -1368 -1399
rect -1302 -1365 -1190 -1359
rect -1302 -1399 -1290 -1365
rect -1202 -1399 -1190 -1365
rect -1302 -1405 -1190 -1399
rect -1124 -1365 -1012 -1359
rect -1124 -1399 -1112 -1365
rect -1024 -1399 -1012 -1365
rect -1124 -1405 -1012 -1399
rect -946 -1365 -834 -1359
rect -946 -1399 -934 -1365
rect -846 -1399 -834 -1365
rect -946 -1405 -834 -1399
rect -768 -1365 -656 -1359
rect -768 -1399 -756 -1365
rect -668 -1399 -656 -1365
rect -768 -1405 -656 -1399
rect -590 -1365 -478 -1359
rect -590 -1399 -578 -1365
rect -490 -1399 -478 -1365
rect -590 -1405 -478 -1399
rect -412 -1365 -300 -1359
rect -412 -1399 -400 -1365
rect -312 -1399 -300 -1365
rect -412 -1405 -300 -1399
rect -234 -1365 -122 -1359
rect -234 -1399 -222 -1365
rect -134 -1399 -122 -1365
rect -234 -1405 -122 -1399
rect -56 -1365 56 -1359
rect -56 -1399 -44 -1365
rect 44 -1399 56 -1365
rect -56 -1405 56 -1399
rect 122 -1365 234 -1359
rect 122 -1399 134 -1365
rect 222 -1399 234 -1365
rect 122 -1405 234 -1399
rect 300 -1365 412 -1359
rect 300 -1399 312 -1365
rect 400 -1399 412 -1365
rect 300 -1405 412 -1399
rect 478 -1365 590 -1359
rect 478 -1399 490 -1365
rect 578 -1399 590 -1365
rect 478 -1405 590 -1399
rect 656 -1365 768 -1359
rect 656 -1399 668 -1365
rect 756 -1399 768 -1365
rect 656 -1405 768 -1399
rect 834 -1365 946 -1359
rect 834 -1399 846 -1365
rect 934 -1399 946 -1365
rect 834 -1405 946 -1399
rect 1012 -1365 1124 -1359
rect 1012 -1399 1024 -1365
rect 1112 -1399 1124 -1365
rect 1012 -1405 1124 -1399
rect 1190 -1365 1302 -1359
rect 1190 -1399 1202 -1365
rect 1290 -1399 1302 -1365
rect 1190 -1405 1302 -1399
rect 1368 -1365 1480 -1359
rect 1368 -1399 1380 -1365
rect 1468 -1399 1480 -1365
rect 1368 -1405 1480 -1399
rect 1546 -1365 1658 -1359
rect 1546 -1399 1558 -1365
rect 1646 -1399 1658 -1365
rect 1546 -1405 1658 -1399
rect 1724 -1365 1836 -1359
rect 1724 -1399 1736 -1365
rect 1824 -1399 1836 -1365
rect 1724 -1405 1836 -1399
rect 1902 -1365 2014 -1359
rect 1902 -1399 1914 -1365
rect 2002 -1399 2014 -1365
rect 1902 -1405 2014 -1399
rect 2080 -1365 2192 -1359
rect 2080 -1399 2092 -1365
rect 2180 -1399 2192 -1365
rect 2080 -1405 2192 -1399
rect 2258 -1365 2370 -1359
rect 2258 -1399 2270 -1365
rect 2358 -1399 2370 -1365
rect 2258 -1405 2370 -1399
rect 2436 -1365 2548 -1359
rect 2436 -1399 2448 -1365
rect 2536 -1399 2548 -1365
rect 2436 -1405 2548 -1399
rect 2614 -1365 2726 -1359
rect 2614 -1399 2626 -1365
rect 2714 -1399 2726 -1365
rect 2614 -1405 2726 -1399
rect 2792 -1365 2904 -1359
rect 2792 -1399 2804 -1365
rect 2892 -1399 2904 -1365
rect 2792 -1405 2904 -1399
rect 2970 -1365 3082 -1359
rect 2970 -1399 2982 -1365
rect 3070 -1399 3082 -1365
rect 2970 -1405 3082 -1399
rect 3148 -1365 3260 -1359
rect 3148 -1399 3160 -1365
rect 3248 -1399 3260 -1365
rect 3148 -1405 3260 -1399
rect 3326 -1365 3438 -1359
rect 3326 -1399 3338 -1365
rect 3426 -1399 3438 -1365
rect 3326 -1405 3438 -1399
rect 3504 -1365 3616 -1359
rect 3504 -1399 3516 -1365
rect 3604 -1399 3616 -1365
rect 3504 -1405 3616 -1399
rect 3682 -1365 3794 -1359
rect 3682 -1399 3694 -1365
rect 3782 -1399 3794 -1365
rect 3682 -1405 3794 -1399
rect 3860 -1365 3972 -1359
rect 3860 -1399 3872 -1365
rect 3960 -1399 3972 -1365
rect 3860 -1405 3972 -1399
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -4119 -1484 4119 1484
string parameters w 6 l 0.6 m 2 nf 45 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
