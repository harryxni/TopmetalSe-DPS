magic
tech sky130A
magscale 1 2
timestamp 1661897893
<< pwell >>
rect -66 -96 366 156
<< nmos >>
rect 20 -70 50 130
rect 250 -70 280 130
<< ndiff >>
rect -40 81 20 130
rect -40 47 -30 81
rect 4 47 20 81
rect -40 13 20 47
rect -40 -21 -30 13
rect 4 -21 20 13
rect -40 -70 20 -21
rect 50 81 120 130
rect 50 47 73 81
rect 107 47 120 81
rect 50 13 120 47
rect 50 -21 73 13
rect 107 -21 120 13
rect 50 -70 120 -21
rect 180 81 250 130
rect 180 47 193 81
rect 227 47 250 81
rect 180 13 250 47
rect 180 -21 193 13
rect 227 -21 250 13
rect 180 -70 250 -21
rect 280 81 340 130
rect 280 47 296 81
rect 330 47 340 81
rect 280 13 340 47
rect 280 -21 296 13
rect 330 -21 340 13
rect 280 -70 340 -21
<< ndiffc >>
rect -30 47 4 81
rect -30 -21 4 13
rect 73 47 107 81
rect 73 -21 107 13
rect 193 47 227 81
rect 193 -21 227 13
rect 296 47 330 81
rect 296 -21 330 13
<< poly >>
rect 238 207 292 223
rect 238 173 248 207
rect 282 173 292 207
rect 20 130 50 160
rect 238 157 292 173
rect 250 130 280 157
rect 20 -100 50 -70
rect 250 -100 280 -70
<< polycont >>
rect 248 173 282 207
<< locali >>
rect 70 207 300 210
rect 70 173 248 207
rect 282 173 300 207
rect 70 170 300 173
rect 70 130 110 170
rect -40 81 4 130
rect -40 47 -30 81
rect -40 13 4 47
rect -40 -21 -30 13
rect -40 -70 4 -21
rect 66 81 110 130
rect 66 47 73 81
rect 107 47 110 81
rect 66 13 110 47
rect 66 -21 73 13
rect 107 -21 110 13
rect 66 -70 110 -21
rect 190 81 234 130
rect 190 47 193 81
rect 227 47 234 81
rect 190 13 234 47
rect 190 -21 193 13
rect 227 -21 234 13
rect 190 -70 234 -21
rect 296 81 340 130
rect 330 47 340 81
rect 296 13 340 47
rect 330 -21 340 13
rect 296 -70 340 -21
rect 190 -80 230 -70
<< labels >>
rlabel locali s 132 186 132 186 4 storage
port 1 nsew
rlabel poly s 33 154 33 154 4 WWL
port 2 nsew
rlabel locali s -37 119 -37 119 4 WBL
port 3 nsew
rlabel locali s 322 -60 322 -60 4 RWL
port 4 nsew
rlabel locali s 216 -74 216 -74 4 RBL
port 5 nsew
<< end >>
