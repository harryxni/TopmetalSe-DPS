magic
tech sky130B
magscale 1 2
timestamp 1662162487
<< locali >>
rect 370 440 410 550
use dram_array  dram_array_0
timestamp 1662162487
transform 1 0 30 0 1 520
box -90 -430 420 370
use dram_array  dram_array_1
timestamp 1662162487
transform 1 0 465 0 1 520
box -90 -430 420 370
<< end >>
