magic
tech sky130B
magscale 1 2
timestamp 1661897893
<< poly >>
rect 60 -65 90 30
rect 60 -323 90 -280
rect 7 -333 90 -323
rect 7 -367 23 -333
rect 57 -365 90 -333
rect 57 -367 73 -365
rect 7 -377 73 -367
<< polycont >>
rect 23 -367 57 -333
<< locali >>
rect 0 307 40 310
rect 0 273 3 307
rect 37 273 40 307
rect 0 210 40 273
rect 350 197 380 230
rect 350 115 380 163
rect 230 20 253 50
rect 0 -123 40 -80
rect 0 -157 3 -123
rect 37 -157 40 -123
rect 0 -160 40 -157
rect 0 -280 40 -260
rect 23 -333 57 -317
rect 23 -383 57 -367
<< viali >>
rect 3 273 37 307
rect 348 163 382 197
rect 253 18 287 52
rect 228 -102 262 -68
rect 3 -157 37 -123
rect 23 -367 57 -333
<< metal1 >>
rect -6 316 46 322
rect -12 264 -6 316
rect 46 264 52 316
rect -6 258 46 264
rect 342 206 388 209
rect 333 154 339 206
rect 391 154 397 206
rect 342 151 388 154
rect 244 61 296 67
rect 244 3 296 9
rect 219 -59 271 -53
rect -10 -114 50 -100
rect 216 -108 219 -62
rect -12 -123 50 -114
rect 271 -108 274 -62
rect 219 -117 271 -111
rect -12 -157 3 -123
rect 37 -157 50 -123
rect -12 -166 50 -157
rect -10 -180 50 -166
rect 78 -180 84 -174
rect -10 -220 84 -180
rect 78 -226 84 -220
rect 136 -226 142 -174
rect 17 -333 63 -321
rect 268 -333 274 -324
rect 17 -367 23 -333
rect 57 -367 274 -333
rect 17 -379 63 -367
rect 268 -376 274 -367
rect 326 -376 332 -324
<< via1 >>
rect -6 307 46 316
rect -6 273 3 307
rect 3 273 37 307
rect 37 273 46 307
rect -6 264 46 273
rect 339 197 391 206
rect 339 163 348 197
rect 348 163 382 197
rect 382 163 391 197
rect 339 154 391 163
rect 244 52 296 61
rect 244 18 253 52
rect 253 18 287 52
rect 287 18 296 52
rect 244 9 296 18
rect 219 -68 271 -59
rect 219 -102 228 -68
rect 228 -102 262 -68
rect 262 -102 271 -68
rect 219 -111 271 -102
rect 84 -226 136 -174
rect 274 -376 326 -324
<< metal2 >>
rect 0 316 40 370
rect -12 264 -6 316
rect 46 264 52 316
rect 0 -430 40 264
rect 175 -50 205 370
rect 339 210 391 212
rect 326 208 404 210
rect 326 152 337 208
rect 393 152 404 208
rect 326 150 404 152
rect 339 148 391 150
rect 261 63 339 65
rect 261 61 272 63
rect 238 9 244 61
rect 261 7 272 9
rect 328 7 339 63
rect 261 5 339 7
rect 175 -59 280 -50
rect 175 -111 219 -59
rect 271 -111 280 -59
rect 175 -120 280 -111
rect 70 -172 140 -160
rect 70 -228 82 -172
rect 138 -228 140 -172
rect 70 -240 140 -228
rect 175 -430 205 -120
rect 274 -320 326 -318
rect 261 -322 339 -320
rect 261 -378 272 -322
rect 328 -378 339 -322
rect 261 -380 339 -378
rect 274 -382 326 -380
<< via2 >>
rect 337 206 393 208
rect 337 154 339 206
rect 339 154 391 206
rect 391 154 393 206
rect 337 152 393 154
rect 272 61 328 63
rect 272 9 296 61
rect 296 9 328 61
rect 272 7 328 9
rect 82 -174 138 -172
rect 82 -226 84 -174
rect 84 -226 136 -174
rect 136 -226 138 -174
rect 82 -228 138 -226
rect 272 -324 328 -322
rect 272 -376 274 -324
rect 274 -376 326 -324
rect 326 -376 328 -324
rect 272 -378 328 -376
<< metal3 >>
rect 330 210 400 215
rect -60 208 420 210
rect -60 152 337 208
rect 393 152 420 208
rect -60 150 420 152
rect 330 145 400 150
rect 265 70 335 76
rect 240 6 268 70
rect 332 6 340 70
rect 240 0 340 6
rect 265 -50 335 0
rect 60 -168 160 -120
rect 60 -232 78 -168
rect 142 -232 160 -168
rect 60 -260 160 -232
rect 265 -320 335 -315
rect -90 -322 420 -320
rect -90 -378 272 -322
rect 328 -378 420 -322
rect -90 -380 420 -378
rect 265 -385 335 -380
<< via3 >>
rect 268 63 332 70
rect 268 7 272 63
rect 272 7 328 63
rect 328 7 332 63
rect 268 6 332 7
rect 78 -172 142 -168
rect 78 -228 82 -172
rect 82 -228 138 -172
rect 138 -228 142 -172
rect 78 -232 142 -228
<< metal4 >>
rect 80 -164 140 370
rect 270 71 330 370
rect 264 70 336 71
rect 264 6 268 70
rect 332 6 336 70
rect 264 5 336 6
rect 74 -168 146 -164
rect 74 -232 78 -168
rect 142 -232 146 -168
rect 74 -236 146 -232
rect 80 -430 140 -236
rect 270 -430 330 5
use dram_cell  dram_cell_0
timestamp 1661897893
transform 1 0 40 0 1 100
box -66 -100 366 223
use dram_cell  dram_cell_1
timestamp 1661897893
transform 1 0 40 0 -1 -150
box -66 -100 366 223
<< end >>
