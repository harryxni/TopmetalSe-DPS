magic
tech sky130B
magscale 1 2
timestamp 1606416512
<< error_p >>
rect -855 372 -797 378
rect -737 372 -679 378
rect -619 372 -561 378
rect -501 372 -443 378
rect -383 372 -325 378
rect -265 372 -207 378
rect -147 372 -89 378
rect -29 372 29 378
rect 89 372 147 378
rect 207 372 265 378
rect 325 372 383 378
rect 443 372 501 378
rect 561 372 619 378
rect 679 372 737 378
rect 797 372 855 378
rect -855 338 -843 372
rect -737 338 -725 372
rect -619 338 -607 372
rect -501 338 -489 372
rect -383 338 -371 372
rect -265 338 -253 372
rect -147 338 -135 372
rect -29 338 -17 372
rect 89 338 101 372
rect 207 338 219 372
rect 325 338 337 372
rect 443 338 455 372
rect 561 338 573 372
rect 679 338 691 372
rect 797 338 809 372
rect -855 332 -797 338
rect -737 332 -679 338
rect -619 332 -561 338
rect -501 332 -443 338
rect -383 332 -325 338
rect -265 332 -207 338
rect -147 332 -89 338
rect -29 332 29 338
rect 89 332 147 338
rect 207 332 265 338
rect 325 332 383 338
rect 443 332 501 338
rect 561 332 619 338
rect 679 332 737 338
rect 797 332 855 338
rect -855 -338 -797 -332
rect -737 -338 -679 -332
rect -619 -338 -561 -332
rect -501 -338 -443 -332
rect -383 -338 -325 -332
rect -265 -338 -207 -332
rect -147 -338 -89 -332
rect -29 -338 29 -332
rect 89 -338 147 -332
rect 207 -338 265 -332
rect 325 -338 383 -332
rect 443 -338 501 -332
rect 561 -338 619 -332
rect 679 -338 737 -332
rect 797 -338 855 -332
rect -855 -372 -843 -338
rect -737 -372 -725 -338
rect -619 -372 -607 -338
rect -501 -372 -489 -338
rect -383 -372 -371 -338
rect -265 -372 -253 -338
rect -147 -372 -135 -338
rect -29 -372 -17 -338
rect 89 -372 101 -338
rect 207 -372 219 -338
rect 325 -372 337 -338
rect 443 -372 455 -338
rect 561 -372 573 -338
rect 679 -372 691 -338
rect 797 -372 809 -338
rect -855 -378 -797 -372
rect -737 -378 -679 -372
rect -619 -378 -561 -372
rect -501 -378 -443 -372
rect -383 -378 -325 -372
rect -265 -378 -207 -372
rect -147 -378 -89 -372
rect -29 -378 29 -372
rect 89 -378 147 -372
rect 207 -378 265 -372
rect 325 -378 383 -372
rect 443 -378 501 -372
rect 561 -378 619 -372
rect 679 -378 737 -372
rect 797 -378 855 -372
<< pwell >>
rect -1052 -510 1052 510
<< nmos >>
rect -856 -300 -796 300
rect -738 -300 -678 300
rect -620 -300 -560 300
rect -502 -300 -442 300
rect -384 -300 -324 300
rect -266 -300 -206 300
rect -148 -300 -88 300
rect -30 -300 30 300
rect 88 -300 148 300
rect 206 -300 266 300
rect 324 -300 384 300
rect 442 -300 502 300
rect 560 -300 620 300
rect 678 -300 738 300
rect 796 -300 856 300
<< ndiff >>
rect -914 288 -856 300
rect -914 -288 -902 288
rect -868 -288 -856 288
rect -914 -300 -856 -288
rect -796 288 -738 300
rect -796 -288 -784 288
rect -750 -288 -738 288
rect -796 -300 -738 -288
rect -678 288 -620 300
rect -678 -288 -666 288
rect -632 -288 -620 288
rect -678 -300 -620 -288
rect -560 288 -502 300
rect -560 -288 -548 288
rect -514 -288 -502 288
rect -560 -300 -502 -288
rect -442 288 -384 300
rect -442 -288 -430 288
rect -396 -288 -384 288
rect -442 -300 -384 -288
rect -324 288 -266 300
rect -324 -288 -312 288
rect -278 -288 -266 288
rect -324 -300 -266 -288
rect -206 288 -148 300
rect -206 -288 -194 288
rect -160 -288 -148 288
rect -206 -300 -148 -288
rect -88 288 -30 300
rect -88 -288 -76 288
rect -42 -288 -30 288
rect -88 -300 -30 -288
rect 30 288 88 300
rect 30 -288 42 288
rect 76 -288 88 288
rect 30 -300 88 -288
rect 148 288 206 300
rect 148 -288 160 288
rect 194 -288 206 288
rect 148 -300 206 -288
rect 266 288 324 300
rect 266 -288 278 288
rect 312 -288 324 288
rect 266 -300 324 -288
rect 384 288 442 300
rect 384 -288 396 288
rect 430 -288 442 288
rect 384 -300 442 -288
rect 502 288 560 300
rect 502 -288 514 288
rect 548 -288 560 288
rect 502 -300 560 -288
rect 620 288 678 300
rect 620 -288 632 288
rect 666 -288 678 288
rect 620 -300 678 -288
rect 738 288 796 300
rect 738 -288 750 288
rect 784 -288 796 288
rect 738 -300 796 -288
rect 856 288 914 300
rect 856 -288 868 288
rect 902 -288 914 288
rect 856 -300 914 -288
<< ndiffc >>
rect -902 -288 -868 288
rect -784 -288 -750 288
rect -666 -288 -632 288
rect -548 -288 -514 288
rect -430 -288 -396 288
rect -312 -288 -278 288
rect -194 -288 -160 288
rect -76 -288 -42 288
rect 42 -288 76 288
rect 160 -288 194 288
rect 278 -288 312 288
rect 396 -288 430 288
rect 514 -288 548 288
rect 632 -288 666 288
rect 750 -288 784 288
rect 868 -288 902 288
<< psubdiff >>
rect -1016 440 -920 474
rect 920 440 1016 474
rect -1016 378 -982 440
rect 982 378 1016 440
rect -1016 -440 -982 -378
rect 982 -440 1016 -378
rect -1016 -474 -920 -440
rect 920 -474 1016 -440
<< psubdiffcont >>
rect -920 440 920 474
rect -1016 -378 -982 378
rect 982 -378 1016 378
rect -920 -474 920 -440
<< poly >>
rect -859 372 -793 388
rect -859 338 -843 372
rect -809 338 -793 372
rect -859 322 -793 338
rect -741 372 -675 388
rect -741 338 -725 372
rect -691 338 -675 372
rect -741 322 -675 338
rect -623 372 -557 388
rect -623 338 -607 372
rect -573 338 -557 372
rect -623 322 -557 338
rect -505 372 -439 388
rect -505 338 -489 372
rect -455 338 -439 372
rect -505 322 -439 338
rect -387 372 -321 388
rect -387 338 -371 372
rect -337 338 -321 372
rect -387 322 -321 338
rect -269 372 -203 388
rect -269 338 -253 372
rect -219 338 -203 372
rect -269 322 -203 338
rect -151 372 -85 388
rect -151 338 -135 372
rect -101 338 -85 372
rect -151 322 -85 338
rect -33 372 33 388
rect -33 338 -17 372
rect 17 338 33 372
rect -33 322 33 338
rect 85 372 151 388
rect 85 338 101 372
rect 135 338 151 372
rect 85 322 151 338
rect 203 372 269 388
rect 203 338 219 372
rect 253 338 269 372
rect 203 322 269 338
rect 321 372 387 388
rect 321 338 337 372
rect 371 338 387 372
rect 321 322 387 338
rect 439 372 505 388
rect 439 338 455 372
rect 489 338 505 372
rect 439 322 505 338
rect 557 372 623 388
rect 557 338 573 372
rect 607 338 623 372
rect 557 322 623 338
rect 675 372 741 388
rect 675 338 691 372
rect 725 338 741 372
rect 675 322 741 338
rect 793 372 859 388
rect 793 338 809 372
rect 843 338 859 372
rect 793 322 859 338
rect -856 300 -796 322
rect -738 300 -678 322
rect -620 300 -560 322
rect -502 300 -442 322
rect -384 300 -324 322
rect -266 300 -206 322
rect -148 300 -88 322
rect -30 300 30 322
rect 88 300 148 322
rect 206 300 266 322
rect 324 300 384 322
rect 442 300 502 322
rect 560 300 620 322
rect 678 300 738 322
rect 796 300 856 322
rect -856 -322 -796 -300
rect -738 -322 -678 -300
rect -620 -322 -560 -300
rect -502 -322 -442 -300
rect -384 -322 -324 -300
rect -266 -322 -206 -300
rect -148 -322 -88 -300
rect -30 -322 30 -300
rect 88 -322 148 -300
rect 206 -322 266 -300
rect 324 -322 384 -300
rect 442 -322 502 -300
rect 560 -322 620 -300
rect 678 -322 738 -300
rect 796 -322 856 -300
rect -859 -338 -793 -322
rect -859 -372 -843 -338
rect -809 -372 -793 -338
rect -859 -388 -793 -372
rect -741 -338 -675 -322
rect -741 -372 -725 -338
rect -691 -372 -675 -338
rect -741 -388 -675 -372
rect -623 -338 -557 -322
rect -623 -372 -607 -338
rect -573 -372 -557 -338
rect -623 -388 -557 -372
rect -505 -338 -439 -322
rect -505 -372 -489 -338
rect -455 -372 -439 -338
rect -505 -388 -439 -372
rect -387 -338 -321 -322
rect -387 -372 -371 -338
rect -337 -372 -321 -338
rect -387 -388 -321 -372
rect -269 -338 -203 -322
rect -269 -372 -253 -338
rect -219 -372 -203 -338
rect -269 -388 -203 -372
rect -151 -338 -85 -322
rect -151 -372 -135 -338
rect -101 -372 -85 -338
rect -151 -388 -85 -372
rect -33 -338 33 -322
rect -33 -372 -17 -338
rect 17 -372 33 -338
rect -33 -388 33 -372
rect 85 -338 151 -322
rect 85 -372 101 -338
rect 135 -372 151 -338
rect 85 -388 151 -372
rect 203 -338 269 -322
rect 203 -372 219 -338
rect 253 -372 269 -338
rect 203 -388 269 -372
rect 321 -338 387 -322
rect 321 -372 337 -338
rect 371 -372 387 -338
rect 321 -388 387 -372
rect 439 -338 505 -322
rect 439 -372 455 -338
rect 489 -372 505 -338
rect 439 -388 505 -372
rect 557 -338 623 -322
rect 557 -372 573 -338
rect 607 -372 623 -338
rect 557 -388 623 -372
rect 675 -338 741 -322
rect 675 -372 691 -338
rect 725 -372 741 -338
rect 675 -388 741 -372
rect 793 -338 859 -322
rect 793 -372 809 -338
rect 843 -372 859 -338
rect 793 -388 859 -372
<< polycont >>
rect -843 338 -809 372
rect -725 338 -691 372
rect -607 338 -573 372
rect -489 338 -455 372
rect -371 338 -337 372
rect -253 338 -219 372
rect -135 338 -101 372
rect -17 338 17 372
rect 101 338 135 372
rect 219 338 253 372
rect 337 338 371 372
rect 455 338 489 372
rect 573 338 607 372
rect 691 338 725 372
rect 809 338 843 372
rect -843 -372 -809 -338
rect -725 -372 -691 -338
rect -607 -372 -573 -338
rect -489 -372 -455 -338
rect -371 -372 -337 -338
rect -253 -372 -219 -338
rect -135 -372 -101 -338
rect -17 -372 17 -338
rect 101 -372 135 -338
rect 219 -372 253 -338
rect 337 -372 371 -338
rect 455 -372 489 -338
rect 573 -372 607 -338
rect 691 -372 725 -338
rect 809 -372 843 -338
<< locali >>
rect -1016 440 -920 474
rect 920 440 1016 474
rect -1016 378 -982 440
rect 982 378 1016 440
rect -859 338 -843 372
rect -809 338 -793 372
rect -741 338 -725 372
rect -691 338 -675 372
rect -623 338 -607 372
rect -573 338 -557 372
rect -505 338 -489 372
rect -455 338 -439 372
rect -387 338 -371 372
rect -337 338 -321 372
rect -269 338 -253 372
rect -219 338 -203 372
rect -151 338 -135 372
rect -101 338 -85 372
rect -33 338 -17 372
rect 17 338 33 372
rect 85 338 101 372
rect 135 338 151 372
rect 203 338 219 372
rect 253 338 269 372
rect 321 338 337 372
rect 371 338 387 372
rect 439 338 455 372
rect 489 338 505 372
rect 557 338 573 372
rect 607 338 623 372
rect 675 338 691 372
rect 725 338 741 372
rect 793 338 809 372
rect 843 338 859 372
rect -902 288 -868 304
rect -902 -304 -868 -288
rect -784 288 -750 304
rect -784 -304 -750 -288
rect -666 288 -632 304
rect -666 -304 -632 -288
rect -548 288 -514 304
rect -548 -304 -514 -288
rect -430 288 -396 304
rect -430 -304 -396 -288
rect -312 288 -278 304
rect -312 -304 -278 -288
rect -194 288 -160 304
rect -194 -304 -160 -288
rect -76 288 -42 304
rect -76 -304 -42 -288
rect 42 288 76 304
rect 42 -304 76 -288
rect 160 288 194 304
rect 160 -304 194 -288
rect 278 288 312 304
rect 278 -304 312 -288
rect 396 288 430 304
rect 396 -304 430 -288
rect 514 288 548 304
rect 514 -304 548 -288
rect 632 288 666 304
rect 632 -304 666 -288
rect 750 288 784 304
rect 750 -304 784 -288
rect 868 288 902 304
rect 868 -304 902 -288
rect -859 -372 -843 -338
rect -809 -372 -793 -338
rect -741 -372 -725 -338
rect -691 -372 -675 -338
rect -623 -372 -607 -338
rect -573 -372 -557 -338
rect -505 -372 -489 -338
rect -455 -372 -439 -338
rect -387 -372 -371 -338
rect -337 -372 -321 -338
rect -269 -372 -253 -338
rect -219 -372 -203 -338
rect -151 -372 -135 -338
rect -101 -372 -85 -338
rect -33 -372 -17 -338
rect 17 -372 33 -338
rect 85 -372 101 -338
rect 135 -372 151 -338
rect 203 -372 219 -338
rect 253 -372 269 -338
rect 321 -372 337 -338
rect 371 -372 387 -338
rect 439 -372 455 -338
rect 489 -372 505 -338
rect 557 -372 573 -338
rect 607 -372 623 -338
rect 675 -372 691 -338
rect 725 -372 741 -338
rect 793 -372 809 -338
rect 843 -372 859 -338
rect -1016 -440 -982 -378
rect 982 -440 1016 -378
rect -1016 -474 -920 -440
rect 920 -474 1016 -440
<< viali >>
rect -843 338 -809 372
rect -725 338 -691 372
rect -607 338 -573 372
rect -489 338 -455 372
rect -371 338 -337 372
rect -253 338 -219 372
rect -135 338 -101 372
rect -17 338 17 372
rect 101 338 135 372
rect 219 338 253 372
rect 337 338 371 372
rect 455 338 489 372
rect 573 338 607 372
rect 691 338 725 372
rect 809 338 843 372
rect -902 -288 -868 288
rect -784 -288 -750 288
rect -666 -288 -632 288
rect -548 -288 -514 288
rect -430 -288 -396 288
rect -312 -288 -278 288
rect -194 -288 -160 288
rect -76 -288 -42 288
rect 42 -288 76 288
rect 160 -288 194 288
rect 278 -288 312 288
rect 396 -288 430 288
rect 514 -288 548 288
rect 632 -288 666 288
rect 750 -288 784 288
rect 868 -288 902 288
rect -843 -372 -809 -338
rect -725 -372 -691 -338
rect -607 -372 -573 -338
rect -489 -372 -455 -338
rect -371 -372 -337 -338
rect -253 -372 -219 -338
rect -135 -372 -101 -338
rect -17 -372 17 -338
rect 101 -372 135 -338
rect 219 -372 253 -338
rect 337 -372 371 -338
rect 455 -372 489 -338
rect 573 -372 607 -338
rect 691 -372 725 -338
rect 809 -372 843 -338
<< metal1 >>
rect -855 372 -797 378
rect -855 338 -843 372
rect -809 338 -797 372
rect -855 332 -797 338
rect -737 372 -679 378
rect -737 338 -725 372
rect -691 338 -679 372
rect -737 332 -679 338
rect -619 372 -561 378
rect -619 338 -607 372
rect -573 338 -561 372
rect -619 332 -561 338
rect -501 372 -443 378
rect -501 338 -489 372
rect -455 338 -443 372
rect -501 332 -443 338
rect -383 372 -325 378
rect -383 338 -371 372
rect -337 338 -325 372
rect -383 332 -325 338
rect -265 372 -207 378
rect -265 338 -253 372
rect -219 338 -207 372
rect -265 332 -207 338
rect -147 372 -89 378
rect -147 338 -135 372
rect -101 338 -89 372
rect -147 332 -89 338
rect -29 372 29 378
rect -29 338 -17 372
rect 17 338 29 372
rect -29 332 29 338
rect 89 372 147 378
rect 89 338 101 372
rect 135 338 147 372
rect 89 332 147 338
rect 207 372 265 378
rect 207 338 219 372
rect 253 338 265 372
rect 207 332 265 338
rect 325 372 383 378
rect 325 338 337 372
rect 371 338 383 372
rect 325 332 383 338
rect 443 372 501 378
rect 443 338 455 372
rect 489 338 501 372
rect 443 332 501 338
rect 561 372 619 378
rect 561 338 573 372
rect 607 338 619 372
rect 561 332 619 338
rect 679 372 737 378
rect 679 338 691 372
rect 725 338 737 372
rect 679 332 737 338
rect 797 372 855 378
rect 797 338 809 372
rect 843 338 855 372
rect 797 332 855 338
rect -908 288 -862 300
rect -908 -288 -902 288
rect -868 -288 -862 288
rect -908 -300 -862 -288
rect -790 288 -744 300
rect -790 -288 -784 288
rect -750 -288 -744 288
rect -790 -300 -744 -288
rect -672 288 -626 300
rect -672 -288 -666 288
rect -632 -288 -626 288
rect -672 -300 -626 -288
rect -554 288 -508 300
rect -554 -288 -548 288
rect -514 -288 -508 288
rect -554 -300 -508 -288
rect -436 288 -390 300
rect -436 -288 -430 288
rect -396 -288 -390 288
rect -436 -300 -390 -288
rect -318 288 -272 300
rect -318 -288 -312 288
rect -278 -288 -272 288
rect -318 -300 -272 -288
rect -200 288 -154 300
rect -200 -288 -194 288
rect -160 -288 -154 288
rect -200 -300 -154 -288
rect -82 288 -36 300
rect -82 -288 -76 288
rect -42 -288 -36 288
rect -82 -300 -36 -288
rect 36 288 82 300
rect 36 -288 42 288
rect 76 -288 82 288
rect 36 -300 82 -288
rect 154 288 200 300
rect 154 -288 160 288
rect 194 -288 200 288
rect 154 -300 200 -288
rect 272 288 318 300
rect 272 -288 278 288
rect 312 -288 318 288
rect 272 -300 318 -288
rect 390 288 436 300
rect 390 -288 396 288
rect 430 -288 436 288
rect 390 -300 436 -288
rect 508 288 554 300
rect 508 -288 514 288
rect 548 -288 554 288
rect 508 -300 554 -288
rect 626 288 672 300
rect 626 -288 632 288
rect 666 -288 672 288
rect 626 -300 672 -288
rect 744 288 790 300
rect 744 -288 750 288
rect 784 -288 790 288
rect 744 -300 790 -288
rect 862 288 908 300
rect 862 -288 868 288
rect 902 -288 908 288
rect 862 -300 908 -288
rect -855 -338 -797 -332
rect -855 -372 -843 -338
rect -809 -372 -797 -338
rect -855 -378 -797 -372
rect -737 -338 -679 -332
rect -737 -372 -725 -338
rect -691 -372 -679 -338
rect -737 -378 -679 -372
rect -619 -338 -561 -332
rect -619 -372 -607 -338
rect -573 -372 -561 -338
rect -619 -378 -561 -372
rect -501 -338 -443 -332
rect -501 -372 -489 -338
rect -455 -372 -443 -338
rect -501 -378 -443 -372
rect -383 -338 -325 -332
rect -383 -372 -371 -338
rect -337 -372 -325 -338
rect -383 -378 -325 -372
rect -265 -338 -207 -332
rect -265 -372 -253 -338
rect -219 -372 -207 -338
rect -265 -378 -207 -372
rect -147 -338 -89 -332
rect -147 -372 -135 -338
rect -101 -372 -89 -338
rect -147 -378 -89 -372
rect -29 -338 29 -332
rect -29 -372 -17 -338
rect 17 -372 29 -338
rect -29 -378 29 -372
rect 89 -338 147 -332
rect 89 -372 101 -338
rect 135 -372 147 -338
rect 89 -378 147 -372
rect 207 -338 265 -332
rect 207 -372 219 -338
rect 253 -372 265 -338
rect 207 -378 265 -372
rect 325 -338 383 -332
rect 325 -372 337 -338
rect 371 -372 383 -338
rect 325 -378 383 -372
rect 443 -338 501 -332
rect 443 -372 455 -338
rect 489 -372 501 -338
rect 443 -378 501 -372
rect 561 -338 619 -332
rect 561 -372 573 -338
rect 607 -372 619 -338
rect 561 -378 619 -372
rect 679 -338 737 -332
rect 679 -372 691 -338
rect 725 -372 737 -338
rect 679 -378 737 -372
rect 797 -338 855 -332
rect 797 -372 809 -338
rect 843 -372 855 -338
rect 797 -378 855 -372
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -999 -457 999 457
string parameters w 3 l 0.3 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
