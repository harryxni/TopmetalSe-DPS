magic
tech sky130A
magscale 1 2
timestamp 1662070103
<< error_s >>
rect 6185 10704 6359 10798
rect 6439 10524 6613 10704
rect 6029 10488 6649 10524
rect 6084 10483 6154 10488
rect 6439 10464 6613 10488
rect 6089 10428 6709 10464
rect 6089 10423 6214 10428
rect 6089 10404 6709 10408
rect 6029 10344 6649 10348
rect 6029 10288 6649 10324
rect 6089 10228 6709 10264
rect 6029 9988 6609 10024
rect 6194 9983 6274 9988
rect 6089 9928 6669 9964
rect 6126 9923 6334 9928
rect 6126 9904 6199 9923
rect 6186 9844 6199 9881
rect 6129 9668 6649 9704
rect 6129 9663 6184 9668
rect 6189 9608 6709 9644
rect 6189 9603 6244 9608
rect 6209 9538 6649 9574
rect 6269 9454 6709 9514
rect 6209 9394 6649 9428
rect 6239 9368 6649 9394
rect 6299 9308 6709 9344
rect 6141 9088 6649 9092
rect 6169 9060 6677 9064
rect 6029 8178 6639 8214
rect 6089 8118 6699 8154
rect 6379 7918 6649 7954
rect 6439 7858 6709 7894
use bottom_left_pixel  bottom_left_pixel_0
timestamp 1662070103
transform 1 0 3089 0 1 4490
box -2819 -4490 3950 3640
use left_pixel  left_pixel_0
timestamp 1662068818
transform 1 0 3089 0 1 7498
box -2819 -148 3560 3640
use top_right_pixel  top_right_pixel_0
timestamp 1662070103
transform 1 0 6169 0 1 7414
box -80 -310 6840 4380
<< end >>
