magic
tech sky130B
magscale 1 2
timestamp 1607735006
<< pwell >>
rect -1947 -810 1947 810
<< nmos >>
rect -1751 -600 -1631 600
rect -1573 -600 -1453 600
rect -1395 -600 -1275 600
rect -1217 -600 -1097 600
rect -1039 -600 -919 600
rect -861 -600 -741 600
rect -683 -600 -563 600
rect -505 -600 -385 600
rect -327 -600 -207 600
rect -149 -600 -29 600
rect 29 -600 149 600
rect 207 -600 327 600
rect 385 -600 505 600
rect 563 -600 683 600
rect 741 -600 861 600
rect 919 -600 1039 600
rect 1097 -600 1217 600
rect 1275 -600 1395 600
rect 1453 -600 1573 600
rect 1631 -600 1751 600
<< ndiff >>
rect -1809 588 -1751 600
rect -1809 -588 -1797 588
rect -1763 -588 -1751 588
rect -1809 -600 -1751 -588
rect -1631 588 -1573 600
rect -1631 -588 -1619 588
rect -1585 -588 -1573 588
rect -1631 -600 -1573 -588
rect -1453 588 -1395 600
rect -1453 -588 -1441 588
rect -1407 -588 -1395 588
rect -1453 -600 -1395 -588
rect -1275 588 -1217 600
rect -1275 -588 -1263 588
rect -1229 -588 -1217 588
rect -1275 -600 -1217 -588
rect -1097 588 -1039 600
rect -1097 -588 -1085 588
rect -1051 -588 -1039 588
rect -1097 -600 -1039 -588
rect -919 588 -861 600
rect -919 -588 -907 588
rect -873 -588 -861 588
rect -919 -600 -861 -588
rect -741 588 -683 600
rect -741 -588 -729 588
rect -695 -588 -683 588
rect -741 -600 -683 -588
rect -563 588 -505 600
rect -563 -588 -551 588
rect -517 -588 -505 588
rect -563 -600 -505 -588
rect -385 588 -327 600
rect -385 -588 -373 588
rect -339 -588 -327 588
rect -385 -600 -327 -588
rect -207 588 -149 600
rect -207 -588 -195 588
rect -161 -588 -149 588
rect -207 -600 -149 -588
rect -29 588 29 600
rect -29 -588 -17 588
rect 17 -588 29 588
rect -29 -600 29 -588
rect 149 588 207 600
rect 149 -588 161 588
rect 195 -588 207 588
rect 149 -600 207 -588
rect 327 588 385 600
rect 327 -588 339 588
rect 373 -588 385 588
rect 327 -600 385 -588
rect 505 588 563 600
rect 505 -588 517 588
rect 551 -588 563 588
rect 505 -600 563 -588
rect 683 588 741 600
rect 683 -588 695 588
rect 729 -588 741 588
rect 683 -600 741 -588
rect 861 588 919 600
rect 861 -588 873 588
rect 907 -588 919 588
rect 861 -600 919 -588
rect 1039 588 1097 600
rect 1039 -588 1051 588
rect 1085 -588 1097 588
rect 1039 -600 1097 -588
rect 1217 588 1275 600
rect 1217 -588 1229 588
rect 1263 -588 1275 588
rect 1217 -600 1275 -588
rect 1395 588 1453 600
rect 1395 -588 1407 588
rect 1441 -588 1453 588
rect 1395 -600 1453 -588
rect 1573 588 1631 600
rect 1573 -588 1585 588
rect 1619 -588 1631 588
rect 1573 -600 1631 -588
rect 1751 588 1809 600
rect 1751 -588 1763 588
rect 1797 -588 1809 588
rect 1751 -600 1809 -588
<< ndiffc >>
rect -1797 -588 -1763 588
rect -1619 -588 -1585 588
rect -1441 -588 -1407 588
rect -1263 -588 -1229 588
rect -1085 -588 -1051 588
rect -907 -588 -873 588
rect -729 -588 -695 588
rect -551 -588 -517 588
rect -373 -588 -339 588
rect -195 -588 -161 588
rect -17 -588 17 588
rect 161 -588 195 588
rect 339 -588 373 588
rect 517 -588 551 588
rect 695 -588 729 588
rect 873 -588 907 588
rect 1051 -588 1085 588
rect 1229 -588 1263 588
rect 1407 -588 1441 588
rect 1585 -588 1619 588
rect 1763 -588 1797 588
<< psubdiff >>
rect -1911 740 -1815 774
rect 1815 740 1911 774
rect -1911 678 -1877 740
rect 1877 678 1911 740
rect -1911 -740 -1877 -678
rect 1877 -740 1911 -678
rect -1911 -774 -1815 -740
rect 1815 -774 1911 -740
<< psubdiffcont >>
rect -1815 740 1815 774
rect -1911 -678 -1877 678
rect 1877 -678 1911 678
rect -1815 -774 1815 -740
<< poly >>
rect -1751 672 -1631 688
rect -1751 638 -1735 672
rect -1647 638 -1631 672
rect -1751 600 -1631 638
rect -1573 672 -1453 688
rect -1573 638 -1557 672
rect -1469 638 -1453 672
rect -1573 600 -1453 638
rect -1395 672 -1275 688
rect -1395 638 -1379 672
rect -1291 638 -1275 672
rect -1395 600 -1275 638
rect -1217 672 -1097 688
rect -1217 638 -1201 672
rect -1113 638 -1097 672
rect -1217 600 -1097 638
rect -1039 672 -919 688
rect -1039 638 -1023 672
rect -935 638 -919 672
rect -1039 600 -919 638
rect -861 672 -741 688
rect -861 638 -845 672
rect -757 638 -741 672
rect -861 600 -741 638
rect -683 672 -563 688
rect -683 638 -667 672
rect -579 638 -563 672
rect -683 600 -563 638
rect -505 672 -385 688
rect -505 638 -489 672
rect -401 638 -385 672
rect -505 600 -385 638
rect -327 672 -207 688
rect -327 638 -311 672
rect -223 638 -207 672
rect -327 600 -207 638
rect -149 672 -29 688
rect -149 638 -133 672
rect -45 638 -29 672
rect -149 600 -29 638
rect 29 672 149 688
rect 29 638 45 672
rect 133 638 149 672
rect 29 600 149 638
rect 207 672 327 688
rect 207 638 223 672
rect 311 638 327 672
rect 207 600 327 638
rect 385 672 505 688
rect 385 638 401 672
rect 489 638 505 672
rect 385 600 505 638
rect 563 672 683 688
rect 563 638 579 672
rect 667 638 683 672
rect 563 600 683 638
rect 741 672 861 688
rect 741 638 757 672
rect 845 638 861 672
rect 741 600 861 638
rect 919 672 1039 688
rect 919 638 935 672
rect 1023 638 1039 672
rect 919 600 1039 638
rect 1097 672 1217 688
rect 1097 638 1113 672
rect 1201 638 1217 672
rect 1097 600 1217 638
rect 1275 672 1395 688
rect 1275 638 1291 672
rect 1379 638 1395 672
rect 1275 600 1395 638
rect 1453 672 1573 688
rect 1453 638 1469 672
rect 1557 638 1573 672
rect 1453 600 1573 638
rect 1631 672 1751 688
rect 1631 638 1647 672
rect 1735 638 1751 672
rect 1631 600 1751 638
rect -1751 -638 -1631 -600
rect -1751 -672 -1735 -638
rect -1647 -672 -1631 -638
rect -1751 -688 -1631 -672
rect -1573 -638 -1453 -600
rect -1573 -672 -1557 -638
rect -1469 -672 -1453 -638
rect -1573 -688 -1453 -672
rect -1395 -638 -1275 -600
rect -1395 -672 -1379 -638
rect -1291 -672 -1275 -638
rect -1395 -688 -1275 -672
rect -1217 -638 -1097 -600
rect -1217 -672 -1201 -638
rect -1113 -672 -1097 -638
rect -1217 -688 -1097 -672
rect -1039 -638 -919 -600
rect -1039 -672 -1023 -638
rect -935 -672 -919 -638
rect -1039 -688 -919 -672
rect -861 -638 -741 -600
rect -861 -672 -845 -638
rect -757 -672 -741 -638
rect -861 -688 -741 -672
rect -683 -638 -563 -600
rect -683 -672 -667 -638
rect -579 -672 -563 -638
rect -683 -688 -563 -672
rect -505 -638 -385 -600
rect -505 -672 -489 -638
rect -401 -672 -385 -638
rect -505 -688 -385 -672
rect -327 -638 -207 -600
rect -327 -672 -311 -638
rect -223 -672 -207 -638
rect -327 -688 -207 -672
rect -149 -638 -29 -600
rect -149 -672 -133 -638
rect -45 -672 -29 -638
rect -149 -688 -29 -672
rect 29 -638 149 -600
rect 29 -672 45 -638
rect 133 -672 149 -638
rect 29 -688 149 -672
rect 207 -638 327 -600
rect 207 -672 223 -638
rect 311 -672 327 -638
rect 207 -688 327 -672
rect 385 -638 505 -600
rect 385 -672 401 -638
rect 489 -672 505 -638
rect 385 -688 505 -672
rect 563 -638 683 -600
rect 563 -672 579 -638
rect 667 -672 683 -638
rect 563 -688 683 -672
rect 741 -638 861 -600
rect 741 -672 757 -638
rect 845 -672 861 -638
rect 741 -688 861 -672
rect 919 -638 1039 -600
rect 919 -672 935 -638
rect 1023 -672 1039 -638
rect 919 -688 1039 -672
rect 1097 -638 1217 -600
rect 1097 -672 1113 -638
rect 1201 -672 1217 -638
rect 1097 -688 1217 -672
rect 1275 -638 1395 -600
rect 1275 -672 1291 -638
rect 1379 -672 1395 -638
rect 1275 -688 1395 -672
rect 1453 -638 1573 -600
rect 1453 -672 1469 -638
rect 1557 -672 1573 -638
rect 1453 -688 1573 -672
rect 1631 -638 1751 -600
rect 1631 -672 1647 -638
rect 1735 -672 1751 -638
rect 1631 -688 1751 -672
<< polycont >>
rect -1735 638 -1647 672
rect -1557 638 -1469 672
rect -1379 638 -1291 672
rect -1201 638 -1113 672
rect -1023 638 -935 672
rect -845 638 -757 672
rect -667 638 -579 672
rect -489 638 -401 672
rect -311 638 -223 672
rect -133 638 -45 672
rect 45 638 133 672
rect 223 638 311 672
rect 401 638 489 672
rect 579 638 667 672
rect 757 638 845 672
rect 935 638 1023 672
rect 1113 638 1201 672
rect 1291 638 1379 672
rect 1469 638 1557 672
rect 1647 638 1735 672
rect -1735 -672 -1647 -638
rect -1557 -672 -1469 -638
rect -1379 -672 -1291 -638
rect -1201 -672 -1113 -638
rect -1023 -672 -935 -638
rect -845 -672 -757 -638
rect -667 -672 -579 -638
rect -489 -672 -401 -638
rect -311 -672 -223 -638
rect -133 -672 -45 -638
rect 45 -672 133 -638
rect 223 -672 311 -638
rect 401 -672 489 -638
rect 579 -672 667 -638
rect 757 -672 845 -638
rect 935 -672 1023 -638
rect 1113 -672 1201 -638
rect 1291 -672 1379 -638
rect 1469 -672 1557 -638
rect 1647 -672 1735 -638
<< locali >>
rect -1911 740 -1815 774
rect 1815 740 1911 774
rect -1911 678 -1877 740
rect 1877 678 1911 740
rect -1751 638 -1735 672
rect -1647 638 -1631 672
rect -1573 638 -1557 672
rect -1469 638 -1453 672
rect -1395 638 -1379 672
rect -1291 638 -1275 672
rect -1217 638 -1201 672
rect -1113 638 -1097 672
rect -1039 638 -1023 672
rect -935 638 -919 672
rect -861 638 -845 672
rect -757 638 -741 672
rect -683 638 -667 672
rect -579 638 -563 672
rect -505 638 -489 672
rect -401 638 -385 672
rect -327 638 -311 672
rect -223 638 -207 672
rect -149 638 -133 672
rect -45 638 -29 672
rect 29 638 45 672
rect 133 638 149 672
rect 207 638 223 672
rect 311 638 327 672
rect 385 638 401 672
rect 489 638 505 672
rect 563 638 579 672
rect 667 638 683 672
rect 741 638 757 672
rect 845 638 861 672
rect 919 638 935 672
rect 1023 638 1039 672
rect 1097 638 1113 672
rect 1201 638 1217 672
rect 1275 638 1291 672
rect 1379 638 1395 672
rect 1453 638 1469 672
rect 1557 638 1573 672
rect 1631 638 1647 672
rect 1735 638 1751 672
rect -1797 588 -1763 604
rect -1797 -604 -1763 -588
rect -1619 588 -1585 604
rect -1619 -604 -1585 -588
rect -1441 588 -1407 604
rect -1441 -604 -1407 -588
rect -1263 588 -1229 604
rect -1263 -604 -1229 -588
rect -1085 588 -1051 604
rect -1085 -604 -1051 -588
rect -907 588 -873 604
rect -907 -604 -873 -588
rect -729 588 -695 604
rect -729 -604 -695 -588
rect -551 588 -517 604
rect -551 -604 -517 -588
rect -373 588 -339 604
rect -373 -604 -339 -588
rect -195 588 -161 604
rect -195 -604 -161 -588
rect -17 588 17 604
rect -17 -604 17 -588
rect 161 588 195 604
rect 161 -604 195 -588
rect 339 588 373 604
rect 339 -604 373 -588
rect 517 588 551 604
rect 517 -604 551 -588
rect 695 588 729 604
rect 695 -604 729 -588
rect 873 588 907 604
rect 873 -604 907 -588
rect 1051 588 1085 604
rect 1051 -604 1085 -588
rect 1229 588 1263 604
rect 1229 -604 1263 -588
rect 1407 588 1441 604
rect 1407 -604 1441 -588
rect 1585 588 1619 604
rect 1585 -604 1619 -588
rect 1763 588 1797 604
rect 1763 -604 1797 -588
rect -1751 -672 -1735 -638
rect -1647 -672 -1631 -638
rect -1573 -672 -1557 -638
rect -1469 -672 -1453 -638
rect -1395 -672 -1379 -638
rect -1291 -672 -1275 -638
rect -1217 -672 -1201 -638
rect -1113 -672 -1097 -638
rect -1039 -672 -1023 -638
rect -935 -672 -919 -638
rect -861 -672 -845 -638
rect -757 -672 -741 -638
rect -683 -672 -667 -638
rect -579 -672 -563 -638
rect -505 -672 -489 -638
rect -401 -672 -385 -638
rect -327 -672 -311 -638
rect -223 -672 -207 -638
rect -149 -672 -133 -638
rect -45 -672 -29 -638
rect 29 -672 45 -638
rect 133 -672 149 -638
rect 207 -672 223 -638
rect 311 -672 327 -638
rect 385 -672 401 -638
rect 489 -672 505 -638
rect 563 -672 579 -638
rect 667 -672 683 -638
rect 741 -672 757 -638
rect 845 -672 861 -638
rect 919 -672 935 -638
rect 1023 -672 1039 -638
rect 1097 -672 1113 -638
rect 1201 -672 1217 -638
rect 1275 -672 1291 -638
rect 1379 -672 1395 -638
rect 1453 -672 1469 -638
rect 1557 -672 1573 -638
rect 1631 -672 1647 -638
rect 1735 -672 1751 -638
rect -1911 -740 -1877 -678
rect 1877 -740 1911 -678
rect -1911 -774 -1815 -740
rect 1815 -774 1911 -740
<< viali >>
rect -1735 638 -1647 672
rect -1557 638 -1469 672
rect -1379 638 -1291 672
rect -1201 638 -1113 672
rect -1023 638 -935 672
rect -845 638 -757 672
rect -667 638 -579 672
rect -489 638 -401 672
rect -311 638 -223 672
rect -133 638 -45 672
rect 45 638 133 672
rect 223 638 311 672
rect 401 638 489 672
rect 579 638 667 672
rect 757 638 845 672
rect 935 638 1023 672
rect 1113 638 1201 672
rect 1291 638 1379 672
rect 1469 638 1557 672
rect 1647 638 1735 672
rect -1797 -588 -1763 588
rect -1619 -588 -1585 588
rect -1441 -588 -1407 588
rect -1263 -588 -1229 588
rect -1085 -588 -1051 588
rect -907 -588 -873 588
rect -729 -588 -695 588
rect -551 -588 -517 588
rect -373 -588 -339 588
rect -195 -588 -161 588
rect -17 -588 17 588
rect 161 -588 195 588
rect 339 -588 373 588
rect 517 -588 551 588
rect 695 -588 729 588
rect 873 -588 907 588
rect 1051 -588 1085 588
rect 1229 -588 1263 588
rect 1407 -588 1441 588
rect 1585 -588 1619 588
rect 1763 -588 1797 588
rect -1735 -672 -1647 -638
rect -1557 -672 -1469 -638
rect -1379 -672 -1291 -638
rect -1201 -672 -1113 -638
rect -1023 -672 -935 -638
rect -845 -672 -757 -638
rect -667 -672 -579 -638
rect -489 -672 -401 -638
rect -311 -672 -223 -638
rect -133 -672 -45 -638
rect 45 -672 133 -638
rect 223 -672 311 -638
rect 401 -672 489 -638
rect 579 -672 667 -638
rect 757 -672 845 -638
rect 935 -672 1023 -638
rect 1113 -672 1201 -638
rect 1291 -672 1379 -638
rect 1469 -672 1557 -638
rect 1647 -672 1735 -638
<< metal1 >>
rect -1747 672 -1635 678
rect -1747 638 -1735 672
rect -1647 638 -1635 672
rect -1747 632 -1635 638
rect -1569 672 -1457 678
rect -1569 638 -1557 672
rect -1469 638 -1457 672
rect -1569 632 -1457 638
rect -1391 672 -1279 678
rect -1391 638 -1379 672
rect -1291 638 -1279 672
rect -1391 632 -1279 638
rect -1213 672 -1101 678
rect -1213 638 -1201 672
rect -1113 638 -1101 672
rect -1213 632 -1101 638
rect -1035 672 -923 678
rect -1035 638 -1023 672
rect -935 638 -923 672
rect -1035 632 -923 638
rect -857 672 -745 678
rect -857 638 -845 672
rect -757 638 -745 672
rect -857 632 -745 638
rect -679 672 -567 678
rect -679 638 -667 672
rect -579 638 -567 672
rect -679 632 -567 638
rect -501 672 -389 678
rect -501 638 -489 672
rect -401 638 -389 672
rect -501 632 -389 638
rect -323 672 -211 678
rect -323 638 -311 672
rect -223 638 -211 672
rect -323 632 -211 638
rect -145 672 -33 678
rect -145 638 -133 672
rect -45 638 -33 672
rect -145 632 -33 638
rect 33 672 145 678
rect 33 638 45 672
rect 133 638 145 672
rect 33 632 145 638
rect 211 672 323 678
rect 211 638 223 672
rect 311 638 323 672
rect 211 632 323 638
rect 389 672 501 678
rect 389 638 401 672
rect 489 638 501 672
rect 389 632 501 638
rect 567 672 679 678
rect 567 638 579 672
rect 667 638 679 672
rect 567 632 679 638
rect 745 672 857 678
rect 745 638 757 672
rect 845 638 857 672
rect 745 632 857 638
rect 923 672 1035 678
rect 923 638 935 672
rect 1023 638 1035 672
rect 923 632 1035 638
rect 1101 672 1213 678
rect 1101 638 1113 672
rect 1201 638 1213 672
rect 1101 632 1213 638
rect 1279 672 1391 678
rect 1279 638 1291 672
rect 1379 638 1391 672
rect 1279 632 1391 638
rect 1457 672 1569 678
rect 1457 638 1469 672
rect 1557 638 1569 672
rect 1457 632 1569 638
rect 1635 672 1747 678
rect 1635 638 1647 672
rect 1735 638 1747 672
rect 1635 632 1747 638
rect -1803 588 -1757 600
rect -1803 -588 -1797 588
rect -1763 -588 -1757 588
rect -1803 -600 -1757 -588
rect -1625 588 -1579 600
rect -1625 -588 -1619 588
rect -1585 -588 -1579 588
rect -1625 -600 -1579 -588
rect -1447 588 -1401 600
rect -1447 -588 -1441 588
rect -1407 -588 -1401 588
rect -1447 -600 -1401 -588
rect -1269 588 -1223 600
rect -1269 -588 -1263 588
rect -1229 -588 -1223 588
rect -1269 -600 -1223 -588
rect -1091 588 -1045 600
rect -1091 -588 -1085 588
rect -1051 -588 -1045 588
rect -1091 -600 -1045 -588
rect -913 588 -867 600
rect -913 -588 -907 588
rect -873 -588 -867 588
rect -913 -600 -867 -588
rect -735 588 -689 600
rect -735 -588 -729 588
rect -695 -588 -689 588
rect -735 -600 -689 -588
rect -557 588 -511 600
rect -557 -588 -551 588
rect -517 -588 -511 588
rect -557 -600 -511 -588
rect -379 588 -333 600
rect -379 -588 -373 588
rect -339 -588 -333 588
rect -379 -600 -333 -588
rect -201 588 -155 600
rect -201 -588 -195 588
rect -161 -588 -155 588
rect -201 -600 -155 -588
rect -23 588 23 600
rect -23 -588 -17 588
rect 17 -588 23 588
rect -23 -600 23 -588
rect 155 588 201 600
rect 155 -588 161 588
rect 195 -588 201 588
rect 155 -600 201 -588
rect 333 588 379 600
rect 333 -588 339 588
rect 373 -588 379 588
rect 333 -600 379 -588
rect 511 588 557 600
rect 511 -588 517 588
rect 551 -588 557 588
rect 511 -600 557 -588
rect 689 588 735 600
rect 689 -588 695 588
rect 729 -588 735 588
rect 689 -600 735 -588
rect 867 588 913 600
rect 867 -588 873 588
rect 907 -588 913 588
rect 867 -600 913 -588
rect 1045 588 1091 600
rect 1045 -588 1051 588
rect 1085 -588 1091 588
rect 1045 -600 1091 -588
rect 1223 588 1269 600
rect 1223 -588 1229 588
rect 1263 -588 1269 588
rect 1223 -600 1269 -588
rect 1401 588 1447 600
rect 1401 -588 1407 588
rect 1441 -588 1447 588
rect 1401 -600 1447 -588
rect 1579 588 1625 600
rect 1579 -588 1585 588
rect 1619 -588 1625 588
rect 1579 -600 1625 -588
rect 1757 588 1803 600
rect 1757 -588 1763 588
rect 1797 -588 1803 588
rect 1757 -600 1803 -588
rect -1747 -638 -1635 -632
rect -1747 -672 -1735 -638
rect -1647 -672 -1635 -638
rect -1747 -678 -1635 -672
rect -1569 -638 -1457 -632
rect -1569 -672 -1557 -638
rect -1469 -672 -1457 -638
rect -1569 -678 -1457 -672
rect -1391 -638 -1279 -632
rect -1391 -672 -1379 -638
rect -1291 -672 -1279 -638
rect -1391 -678 -1279 -672
rect -1213 -638 -1101 -632
rect -1213 -672 -1201 -638
rect -1113 -672 -1101 -638
rect -1213 -678 -1101 -672
rect -1035 -638 -923 -632
rect -1035 -672 -1023 -638
rect -935 -672 -923 -638
rect -1035 -678 -923 -672
rect -857 -638 -745 -632
rect -857 -672 -845 -638
rect -757 -672 -745 -638
rect -857 -678 -745 -672
rect -679 -638 -567 -632
rect -679 -672 -667 -638
rect -579 -672 -567 -638
rect -679 -678 -567 -672
rect -501 -638 -389 -632
rect -501 -672 -489 -638
rect -401 -672 -389 -638
rect -501 -678 -389 -672
rect -323 -638 -211 -632
rect -323 -672 -311 -638
rect -223 -672 -211 -638
rect -323 -678 -211 -672
rect -145 -638 -33 -632
rect -145 -672 -133 -638
rect -45 -672 -33 -638
rect -145 -678 -33 -672
rect 33 -638 145 -632
rect 33 -672 45 -638
rect 133 -672 145 -638
rect 33 -678 145 -672
rect 211 -638 323 -632
rect 211 -672 223 -638
rect 311 -672 323 -638
rect 211 -678 323 -672
rect 389 -638 501 -632
rect 389 -672 401 -638
rect 489 -672 501 -638
rect 389 -678 501 -672
rect 567 -638 679 -632
rect 567 -672 579 -638
rect 667 -672 679 -638
rect 567 -678 679 -672
rect 745 -638 857 -632
rect 745 -672 757 -638
rect 845 -672 857 -638
rect 745 -678 857 -672
rect 923 -638 1035 -632
rect 923 -672 935 -638
rect 1023 -672 1035 -638
rect 923 -678 1035 -672
rect 1101 -638 1213 -632
rect 1101 -672 1113 -638
rect 1201 -672 1213 -638
rect 1101 -678 1213 -672
rect 1279 -638 1391 -632
rect 1279 -672 1291 -638
rect 1379 -672 1391 -638
rect 1279 -678 1391 -672
rect 1457 -638 1569 -632
rect 1457 -672 1469 -638
rect 1557 -672 1569 -638
rect 1457 -678 1569 -672
rect 1635 -638 1747 -632
rect 1635 -672 1647 -638
rect 1735 -672 1747 -638
rect 1635 -678 1747 -672
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1894 -757 1894 757
string parameters w 6 l 0.6 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
