magic
tech sky130B
magscale 1 2
timestamp 1608255150
<< nwell >>
rect -211 -327 211 327
<< pmos >>
rect -15 -108 15 108
<< pdiff >>
rect -73 96 -15 108
rect -73 -96 -61 96
rect -27 -96 -15 96
rect -73 -108 -15 -96
rect 15 96 73 108
rect 15 -96 27 96
rect 61 -96 73 96
rect 15 -108 73 -96
<< pdiffc >>
rect -61 -96 -27 96
rect 27 -96 61 96
<< nsubdiff >>
rect -175 257 -79 291
rect 79 257 175 291
rect -175 195 -141 257
rect 141 195 175 257
rect -175 -238 -141 -195
rect 141 -238 175 -195
<< nsubdiffcont >>
rect -79 257 79 291
rect -175 -195 -141 195
rect 141 -195 175 195
<< poly >>
rect -15 108 15 152
rect -15 -145 15 -108
<< locali >>
rect -175 257 -79 291
rect 79 257 175 291
rect -175 195 -141 257
rect 141 195 175 257
rect -61 96 -27 112
rect -61 -112 -27 -96
rect 27 96 61 112
rect 27 -112 61 -96
rect -175 -238 -141 -195
rect 141 -238 175 -195
<< viali >>
rect -61 -96 -27 96
rect 27 -96 61 96
<< metal1 >>
rect -67 96 -21 108
rect -67 -96 -61 96
rect -27 -96 -21 96
rect -67 -108 -21 -96
rect 21 96 67 108
rect 21 -96 27 96
rect 61 -96 67 96
rect 21 -108 67 -96
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -158 -274 158 274
string parameters w 1.08 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
