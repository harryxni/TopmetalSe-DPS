magic
tech sky130B
magscale 1 2
timestamp 1662155535
<< metal1 >>
rect 24140 692850 26600 692870
rect 22490 692780 26600 692850
rect 22490 691070 22560 692780
rect 26520 691070 26600 692780
rect 22490 690940 26600 691070
rect 24140 690410 26600 690940
rect 26190 689470 39770 689570
rect 26190 688990 36060 689470
rect 26200 687790 36060 688990
rect 39510 689460 39770 689470
rect 39510 687790 42700 689460
rect 26200 687620 42700 687790
rect 26663 683632 27687 687620
rect 29716 683675 30585 687620
rect 31111 683649 31609 687620
rect 36390 686900 42700 687620
rect 31111 683145 31609 683151
rect 29716 682800 30585 682806
rect 26663 682322 27687 682328
rect 53715 205825 59960 206575
rect 44080 204950 46260 205280
rect 53879 204990 53991 205825
rect 54079 204990 54191 205825
rect 54279 204990 54391 205825
rect 54479 204990 54591 205825
rect 54679 204990 54791 205825
rect 54879 204990 54991 205825
rect 55079 204990 55191 205825
rect 55279 204990 55391 205825
rect 55479 204990 55591 205825
rect 55679 204990 55791 205825
rect 59210 204990 59960 205825
rect 545850 205030 549270 205460
rect 60625 204990 549270 205030
rect 44080 201770 44290 204950
rect 46040 203890 46260 204950
rect 53720 204960 549270 204990
rect 53720 204930 60690 204960
rect 53720 204740 55880 204930
rect 57195 204740 60690 204930
rect 53720 204700 60690 204740
rect 49580 204410 49640 204416
rect 49640 204350 53720 204410
rect 49580 204344 49640 204350
rect 53660 204120 53720 204350
rect 53520 203905 53610 204120
rect 53405 203890 53765 203905
rect 46040 203870 53765 203890
rect 53490 203835 53765 203870
rect 53490 203645 53680 203835
rect 53490 203470 53685 203645
rect 46040 203370 53685 203470
rect 46040 203360 53630 203370
rect 46040 203342 53670 203360
rect 46040 203297 53685 203342
rect 46040 203170 53580 203297
rect 56375 203170 57125 204700
rect 58105 203170 58855 204700
rect 59210 203170 59960 204700
rect 60625 203170 60690 204700
rect 46040 202800 46260 203170
rect 52270 202800 52570 203170
rect 46040 202500 52570 202800
rect 56225 202620 60690 203170
rect 46040 202040 46260 202500
rect 52270 202040 52570 202500
rect 55570 202500 60690 202620
rect 548610 202500 549270 204960
rect 55570 202490 60730 202500
rect 55570 202470 59960 202490
rect 55550 202420 59960 202470
rect 46040 201770 52570 202040
rect 44080 201740 52570 201770
rect 44080 201560 46260 201740
rect 52270 201070 52570 201740
rect 44914 200770 44920 201070
rect 45220 200770 52570 201070
rect 52270 200130 52570 200770
rect 45014 199830 45020 200130
rect 45320 199830 52570 200130
rect 52270 199110 52570 199830
rect 56060 201090 56260 202420
rect 56590 201090 56790 202420
rect 56060 200890 56790 201090
rect 56060 199720 56260 200890
rect 57320 199720 57520 202420
rect 56060 199520 57520 199720
rect 56060 199110 56260 199520
rect 58170 199110 58370 202420
rect 545850 202320 549270 202500
rect 45444 198810 45450 199110
rect 45750 198950 52980 199110
rect 45750 198850 53000 198950
rect 45750 198810 52980 198850
rect 53170 196510 53270 198950
rect 53510 196530 53610 198880
rect 53870 196530 53970 198950
rect 53164 196410 53170 196510
rect 53270 196410 53276 196510
rect 53504 196430 53510 196530
rect 53610 196430 53616 196530
rect 53870 196424 53970 196430
rect 54230 196430 54330 198950
rect 54590 196480 54690 198950
rect 54590 196374 54690 196380
rect 54950 196430 55050 198950
rect 54230 196324 54330 196330
rect 54950 196324 55050 196330
rect 55310 196350 55410 198950
rect 56060 198910 58370 199110
rect 56060 198890 56260 198910
rect 55310 196250 55760 196350
rect 55860 196250 55866 196350
<< via1 >>
rect 22560 691070 26520 692780
rect 36060 687790 39510 689470
rect 26663 682328 27687 683632
rect 29716 682806 30585 683675
rect 31111 683151 31609 683649
rect 44290 203870 46040 204950
rect 55880 204740 57195 204930
rect 49580 204350 49640 204410
rect 44290 203470 53490 203870
rect 44290 201770 46040 203470
rect 60690 202500 548610 204960
rect 44920 200770 45220 201070
rect 45020 199830 45320 200130
rect 45450 198810 45750 199110
rect 53170 196410 53270 196510
rect 53510 196430 53610 196530
rect 53870 196430 53970 196530
rect 54230 196330 54330 196430
rect 54590 196380 54690 196480
rect 54950 196330 55050 196430
rect 55760 196250 55860 196350
<< metal2 >>
rect 165590 697195 165599 699685
rect 168089 697195 168098 699685
rect 24140 692850 26600 692870
rect 22490 692780 26600 692850
rect 22490 691070 22560 692780
rect 26520 691070 26600 692780
rect 22490 690940 26600 691070
rect 2500 690175 5000 690600
rect 24140 690410 24300 690940
rect 24830 690410 26600 690940
rect 2500 690080 25285 690175
rect 795 690030 25500 690080
rect 2500 688525 25285 690030
rect 2500 685237 5000 688525
rect 2496 682747 2505 685237
rect 4995 682747 5004 685237
rect 29716 683675 30585 683684
rect 26663 683632 27687 683641
rect 2500 682742 5000 682747
rect 26657 682328 26663 683632
rect 27687 682328 27693 683632
rect 29710 682806 29716 683675
rect 30585 682806 30591 683675
rect 31111 683649 31609 683658
rect 31105 683151 31111 683649
rect 31609 683151 31615 683649
rect 31111 683142 31609 683151
rect 29716 682797 30585 682806
rect 26663 682319 27687 682328
rect 32590 206138 32670 689740
rect 33290 207748 33370 689730
rect 33290 207692 33302 207748
rect 33358 207692 33370 207748
rect 33290 207480 33370 207692
rect 32590 206082 32592 206138
rect 32648 206082 32670 206138
rect 32590 193540 32670 206082
rect 34420 199300 34500 689730
rect 35960 689470 39580 689550
rect 35960 687790 36060 689470
rect 39510 689460 39580 689470
rect 39510 689345 42700 689460
rect 39510 687790 40195 689345
rect 35960 687690 40195 687790
rect 35990 686895 40195 687690
rect 42645 686900 42700 689345
rect 42645 686895 42650 686900
rect 35990 686890 42650 686895
rect 40195 686886 42645 686890
rect 54101 211840 54110 211900
rect 54170 211840 54179 211900
rect 44080 204950 46260 205280
rect 44080 201770 44290 204950
rect 46040 204150 46260 204950
rect 54120 204770 54160 211840
rect 54500 209860 54509 209920
rect 54569 209860 54578 209920
rect 54519 204770 54559 209860
rect 54935 207480 54944 207540
rect 55004 207480 55013 207540
rect 54954 204770 54994 207480
rect 56530 205690 56590 205699
rect 56530 205621 56590 205630
rect 55389 205100 55429 205110
rect 56540 205100 56580 205621
rect 55389 205060 56590 205100
rect 55389 204620 55429 205060
rect 545850 205030 549270 205460
rect 60625 204980 549270 205030
rect 55830 204960 549270 204980
rect 55830 204930 60690 204960
rect 55830 204740 55880 204930
rect 60615 204740 60690 204930
rect 55830 204710 60690 204740
rect 49580 204410 49640 204419
rect 49574 204350 49580 204410
rect 49640 204350 49646 204410
rect 49580 204341 49640 204350
rect 46040 203890 53610 204150
rect 46040 203870 53620 203890
rect 53490 203470 53620 203870
rect 46040 203410 53620 203470
rect 46040 201770 46260 203410
rect 53160 203085 53200 203090
rect 53160 203055 53949 203085
rect 53160 202790 53200 203055
rect 54350 203000 54390 203090
rect 55224 203082 55254 203085
rect 54789 203055 54819 203080
rect 53500 202998 53560 203000
rect 53493 202942 53502 202998
rect 53558 202942 53567 202998
rect 53840 202960 54390 203000
rect 54625 203025 54819 203055
rect 53500 202760 53560 202942
rect 53840 202790 53880 202960
rect 54231 202860 54287 202867
rect 54170 202858 54300 202860
rect 54170 202802 54231 202858
rect 54287 202802 54300 202858
rect 54625 202830 54655 203025
rect 54840 202968 54900 202970
rect 54833 202912 54842 202968
rect 54898 202912 54907 202968
rect 54170 202730 54300 202802
rect 54520 202790 54655 202830
rect 54525 202785 54655 202790
rect 54840 202770 54900 202912
rect 55208 202785 55254 203082
rect 55530 202948 55590 202950
rect 55523 202892 55532 202948
rect 55588 202892 55597 202948
rect 55530 202770 55590 202892
rect 60625 202500 60690 204710
rect 548610 202500 549270 204960
rect 545850 202320 549270 202500
rect 44080 201560 46260 201770
rect 44920 201070 45220 201076
rect 44911 200770 44920 201070
rect 45220 200770 45229 201070
rect 44920 200764 45220 200770
rect 45020 200130 45320 200136
rect 45011 199830 45020 200130
rect 45320 199830 45329 200130
rect 45020 199824 45320 199830
rect 48460 199310 51040 199330
rect 48460 199300 48480 199310
rect 34420 199220 48480 199300
rect 48460 199180 48480 199220
rect 51020 199180 51040 199310
rect 48460 199170 51040 199180
rect 45450 199110 45750 199116
rect 45441 198810 45450 199110
rect 45750 198810 45759 199110
rect 45450 198804 45750 198810
rect 53510 196530 53610 196536
rect 53870 196530 53970 196539
rect 53170 196510 53270 196516
rect 53161 196410 53170 196510
rect 53270 196410 53279 196510
rect 53501 196430 53510 196530
rect 53610 196430 53619 196530
rect 53864 196430 53870 196530
rect 53970 196430 53976 196530
rect 54590 196480 54690 196489
rect 54584 196470 54590 196480
rect 54200 196430 54350 196460
rect 53510 196424 53610 196430
rect 53870 196421 53970 196430
rect 53170 196404 53270 196410
rect 54200 196330 54230 196430
rect 54330 196330 54350 196430
rect 54581 196380 54590 196470
rect 54690 196470 54696 196480
rect 54690 196380 54699 196470
rect 54950 196430 55050 196439
rect 54590 196371 54690 196380
rect 54944 196330 54950 196430
rect 55050 196330 55056 196430
rect 55760 196350 55860 196356
rect 54200 196280 54350 196330
rect 54950 196321 55050 196330
rect 55751 196250 55760 196350
rect 55860 196250 55869 196350
rect 55760 196244 55860 196250
rect 75730 26498 75790 26500
rect 75723 26442 75732 26498
rect 75788 26442 75797 26498
rect 75730 10626 75790 26442
rect 72344 10514 155478 10626
rect 75730 10320 75790 10514
rect 69764 8646 69876 8655
rect 68454 8534 69764 8646
rect 69876 8534 151932 8646
rect 69764 8525 69876 8534
rect 66364 7086 66476 7095
rect 64844 6974 66364 7086
rect 66476 6974 148386 7086
rect 66364 6965 66476 6974
rect 62874 5706 62986 5715
rect 56514 5594 62874 5706
rect 62986 5594 144840 5706
rect 62874 5585 62986 5594
rect 55244 4376 55356 4385
rect 54284 4264 55244 4376
rect 55356 4264 141294 4376
rect 55244 4255 55356 4264
rect 52334 3346 52446 3355
rect 50394 3234 52334 3346
rect 52446 3234 137748 3346
rect 52334 3225 52446 3234
rect 49534 2266 49646 2275
rect 47484 2154 49534 2266
rect 49646 2154 134202 2266
rect 49534 2145 49646 2154
rect 46414 1726 46526 1735
rect 44074 1614 46414 1726
rect 46526 1614 130656 1726
rect 46414 1605 46526 1614
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 1614
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 2154
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 3234
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 4264
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 5594
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 6974
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 8534
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 10514
rect 551336 10576 551448 10936
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 10464
rect 576158 9736 576270 10116
rect 576149 9624 576158 9736
rect 576270 9624 576279 9736
rect 558428 7876 558540 8316
rect 554882 6156 554994 7226
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 6044
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 7764
rect 572612 6556 572724 6686
rect 561974 6076 562086 6356
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 5964
rect 565520 6306 565632 6406
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 6194
rect 569066 6286 569178 6466
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 6174
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 6444
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 9624
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 165599 697195 168089 699685
rect 22560 691070 26520 692780
rect 24300 690410 24830 690940
rect 2505 682747 4995 685237
rect 26663 682328 27687 683632
rect 29716 682806 30585 683675
rect 31111 683151 31609 683649
rect 33302 207692 33358 207748
rect 32592 206082 32648 206138
rect 40195 686895 42645 689345
rect 54110 211840 54170 211900
rect 44290 203870 46040 204950
rect 54509 209860 54569 209920
rect 54944 207480 55004 207540
rect 56530 205630 56590 205690
rect 55880 204740 57195 204930
rect 57195 204740 60615 204930
rect 49580 204350 49640 204410
rect 44290 203470 53490 203870
rect 44290 201770 46040 203470
rect 53502 202942 53558 202998
rect 54231 202802 54287 202858
rect 54842 202912 54898 202968
rect 55532 202892 55588 202948
rect 60690 202500 548610 204960
rect 44920 200770 45220 201070
rect 45020 199830 45320 200130
rect 48480 199180 51020 199310
rect 45450 198810 45750 199110
rect 53170 196410 53270 196510
rect 53510 196430 53610 196530
rect 53870 196430 53970 196530
rect 54230 196330 54330 196430
rect 54590 196380 54690 196480
rect 54950 196330 55050 196430
rect 55760 196250 55860 196350
rect 75732 26442 75788 26498
rect 69764 8534 69876 8646
rect 66364 6974 66476 7086
rect 62874 5594 62986 5706
rect 55244 4264 55356 4376
rect 52334 3234 52446 3346
rect 49534 2154 49646 2266
rect 46414 1614 46526 1726
rect 551336 10464 551448 10576
rect 576158 9624 576270 9736
rect 558428 7764 558540 7876
rect 554882 6044 554994 6156
rect 561974 5964 562086 6076
rect 565520 6194 565632 6306
rect 569066 6174 569178 6286
rect 572612 6444 572724 6556
<< metal3 >>
rect 16194 703310 21194 704800
rect 16194 702300 27065 703310
rect 18694 701630 27065 702300
rect 68194 702300 73194 704800
rect 120194 702740 125194 704800
rect 75620 702300 125194 702740
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702310 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 420980 702300 470394 702310
rect 566594 702300 571594 704800
rect 68194 701860 70694 702300
rect 18694 699900 27220 701630
rect 68140 700540 70694 701860
rect 29770 699960 70694 700540
rect 24590 695880 25050 695886
rect 22584 695320 22590 695780
rect 23050 695320 23056 695780
rect 23590 695770 24050 695776
rect 22590 692850 23050 695320
rect 23590 692850 24050 695310
rect 24590 692870 25050 695420
rect 25590 695880 26050 695886
rect 25590 692870 26050 695420
rect 24140 692850 26600 692870
rect 22490 692780 26600 692850
rect 22490 691070 22560 692780
rect 26520 691070 26600 692780
rect 22490 690940 26600 691070
rect 22490 690410 24300 690940
rect 24830 690410 26600 690940
rect 27020 690560 27220 699900
rect 27530 699760 70694 699960
rect 27530 690590 27730 699760
rect 29770 699360 70694 699760
rect 75620 701700 124910 702300
rect 29770 699320 70270 699360
rect 75620 698120 76660 701700
rect 319171 701179 321669 701185
rect 164800 700260 168840 700320
rect 28410 697080 76660 698120
rect 77320 699689 168890 700260
rect 218481 700130 220979 700135
rect 77320 699240 165595 699689
rect -800 685237 5000 685242
rect -800 682747 2505 685237
rect 4995 682747 5000 685237
rect -800 682742 5000 682747
rect -800 680242 1700 682742
rect 22490 680270 24950 690410
rect 28410 690390 29450 697080
rect 77320 695140 78340 699240
rect 164800 697400 165595 699240
rect 165589 697191 165595 697400
rect 168093 699240 168890 699689
rect 215230 700129 220980 700130
rect 215230 699305 218481 700129
rect 168093 697400 168840 699240
rect 172955 698835 218481 699305
rect 168093 697191 168099 697400
rect 165594 697190 168094 697191
rect 30220 694120 78340 695140
rect 30220 690370 31240 694120
rect 172955 693615 173425 698835
rect 215230 697631 218481 698835
rect 220979 697631 220980 700129
rect 215230 697630 220980 697631
rect 224425 699655 319171 700125
rect 218481 697625 220979 697630
rect 32150 693145 173425 693615
rect 32150 691050 32620 693145
rect 33300 692645 33770 692675
rect 224425 692645 224895 699655
rect 319171 698675 321669 698681
rect 33300 692175 224895 692645
rect 33300 691000 33770 692175
rect 34660 691430 35130 691620
rect 415560 691430 418060 702300
rect 34660 690960 418060 691430
rect 415560 690760 418060 690960
rect 420980 699810 467894 702300
rect 26500 684896 26590 689773
rect 29711 683675 30590 683680
rect 29711 683670 29716 683675
rect 30585 683670 30590 683675
rect 26658 683632 27692 683637
rect 26658 683627 26663 683632
rect 27687 683627 27692 683632
rect 31106 683649 31614 683654
rect 31106 683644 31111 683649
rect 31609 683644 31614 683649
rect 31106 683140 31614 683146
rect 29711 682795 30590 682801
rect 26658 682317 27692 682323
rect 22484 678880 22490 680270
rect 18410 677810 22490 678880
rect 24950 677810 24956 680270
rect 18410 676420 24950 677810
rect 18410 648642 20870 676420
rect -800 646182 20870 648642
rect -800 643842 1660 646182
rect -800 637210 1660 638642
rect -800 634750 19000 637210
rect 21460 634750 21466 637210
rect -800 633842 1660 634750
rect -800 562060 1660 564242
rect -800 559600 14060 562060
rect 16520 559600 16526 562060
rect -800 559442 1660 559600
rect -800 552210 1660 554242
rect -800 549750 14400 552210
rect 16860 549750 16866 552210
rect -800 549442 1660 549750
rect 35680 511660 35880 690760
rect 36240 689349 42840 689740
rect 36240 686891 40191 689349
rect 42649 686891 42840 689349
rect 420980 686930 423480 699810
rect 36240 686560 42840 686891
rect 1360 511642 35880 511660
rect -800 511530 35880 511642
rect 1360 511460 35880 511530
rect 35680 510910 35880 511460
rect 46460 684430 423480 686930
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect -800 295420 36783 295532
rect 36895 295420 36901 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect -800 252398 30075 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect 29941 250039 30053 252398
rect 29941 249971 29956 250039
rect 30024 249971 30053 250039
rect 29941 249942 30053 249971
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect -800 214888 1660 219688
rect 46460 215520 48960 684430
rect 582300 677984 584800 682984
rect 576090 644330 584800 644584
rect 576030 639784 584800 644330
rect 576030 634584 580530 639784
rect 576030 632260 584800 634584
rect 546150 629800 584800 632260
rect 46460 213020 52500 215520
rect -800 204888 1660 209688
rect 33297 207750 33363 207753
rect 33297 207748 50340 207750
rect 33297 207692 33302 207748
rect 33358 207692 50340 207748
rect 33297 207690 50340 207692
rect 33297 207687 33363 207690
rect 32550 206142 32700 206170
rect 32550 206078 32588 206142
rect 32652 206078 32700 206142
rect 32550 206040 32700 206078
rect 43890 204950 46350 205720
rect 43890 204858 44290 204950
rect 24944 203217 24950 204858
rect 26591 203217 44290 204858
rect 46040 204150 46350 204950
rect 49500 204415 49710 204500
rect 49500 204351 49575 204415
rect 49645 204351 49710 204415
rect 50280 204460 50340 207690
rect 51420 204630 51480 213020
rect 54050 211905 54210 211940
rect 54050 211900 54111 211905
rect 54050 211840 54110 211900
rect 54050 211835 54111 211840
rect 54175 211835 54210 211905
rect 54050 211760 54210 211835
rect 54480 209925 54640 209970
rect 54480 209920 54510 209925
rect 54480 209860 54509 209920
rect 54480 209855 54510 209860
rect 54574 209855 54640 209925
rect 54480 209840 54640 209855
rect 54870 207545 55100 207570
rect 54870 207540 54945 207545
rect 54870 207480 54944 207540
rect 54870 207475 54945 207480
rect 55009 207475 55100 207545
rect 54870 207390 55100 207475
rect 546150 206970 548610 629800
rect 582340 629784 584800 629800
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect 56480 205695 56640 205750
rect 56480 205631 56525 205695
rect 56595 205631 56640 205695
rect 56480 205630 56530 205631
rect 56590 205630 56640 205631
rect 56480 205590 56640 205630
rect 546150 205030 549530 206970
rect 60625 204970 549530 205030
rect 53760 204960 549530 204970
rect 53760 204930 60690 204960
rect 53760 204820 55880 204930
rect 53670 204740 55880 204820
rect 60615 204740 60690 204930
rect 53670 204710 60690 204740
rect 53670 204700 55480 204710
rect 51360 204570 55530 204630
rect 50280 204400 55610 204460
rect 49500 204350 49580 204351
rect 49640 204350 49710 204351
rect 49500 204310 49710 204350
rect 46040 203890 53610 204150
rect 46040 203870 53620 203890
rect 53490 203470 53620 203870
rect 43890 201770 44290 203217
rect 46040 203410 53620 203470
rect 46040 201770 46350 203410
rect 51754 203210 53660 203270
rect 51754 203032 51814 203210
rect 51752 203026 51816 203032
rect 51752 202956 51816 202962
rect 53480 203002 53600 203020
rect 53480 202938 53498 203002
rect 53562 202938 53600 203002
rect 53480 202920 53600 202938
rect 54820 202972 54910 202990
rect 54820 202908 54838 202972
rect 54902 202908 54910 202972
rect 54820 202880 54910 202908
rect 55510 202952 55630 202990
rect 55510 202888 55528 202952
rect 55592 202888 55630 202952
rect 55510 202880 55630 202888
rect 54227 202863 54291 202868
rect 54226 202862 54292 202863
rect 54226 202860 54227 202862
rect 54170 202798 54227 202860
rect 54291 202860 54292 202862
rect 54291 202798 54300 202860
rect 54170 202730 54300 202798
rect 60625 202500 60690 204710
rect 548610 202500 549530 204960
rect 43890 201075 46350 201770
rect 59565 201630 549530 202500
rect 547970 201620 549530 201630
rect 24649 200765 25772 200771
rect 43890 200765 44915 201075
rect 45215 201070 46350 201075
rect 45220 200770 46350 201070
rect 45215 200765 46350 200770
rect 24643 199640 24649 200765
rect 25774 200135 46350 200765
rect 25774 199825 45015 200135
rect 45315 200130 46350 200135
rect 45320 199830 46350 200130
rect 45315 199825 46350 199830
rect 25774 199640 46350 199825
rect 24649 199634 25772 199640
rect 43890 199115 46350 199640
rect 49178 199490 49184 199560
rect 49254 199490 52935 199560
rect 48460 199310 51040 199330
rect 48460 199180 48480 199310
rect 51020 199240 51040 199310
rect 51020 199180 52930 199240
rect 48460 199170 51040 199180
rect 43890 198805 45445 199115
rect 45745 199110 46350 199115
rect 45750 198810 46350 199110
rect 45745 198805 46350 198810
rect 24781 197784 27239 197790
rect 43890 197784 46350 198805
rect 24775 195324 24781 197784
rect 27241 196650 46350 197784
rect 27241 196530 57890 196650
rect 27241 196510 53510 196530
rect 27241 196410 53170 196510
rect 53270 196430 53510 196510
rect 53610 196430 53870 196530
rect 53970 196480 57890 196530
rect 53970 196430 54590 196480
rect 53270 196410 54230 196430
rect 27241 196330 54230 196410
rect 54330 196380 54590 196430
rect 54690 196430 57890 196480
rect 54690 196380 54950 196430
rect 54330 196330 54950 196380
rect 55050 196355 57890 196430
rect 55050 196350 55765 196355
rect 55050 196330 55760 196350
rect 27241 196250 55760 196330
rect 27241 196245 55765 196250
rect 55865 196245 57890 196355
rect 27241 195324 57890 196245
rect 24781 195318 27239 195324
rect 43890 194190 57890 195324
rect 24930 191312 27388 191318
rect 43890 191312 46350 194190
rect 582340 191430 584800 196230
rect 24924 188852 24930 191312
rect 27390 188852 46350 191312
rect 24930 188846 27388 188852
rect 43890 184967 46350 188852
rect 24633 182507 24639 184967
rect 27099 182507 46350 184967
rect -800 172888 1660 177688
rect -800 165348 1660 167688
rect 43890 165348 46350 182507
rect 582340 181430 584800 186230
rect -800 162888 3213 165348
rect 39658 162888 46350 165348
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 75680 26502 75850 26540
rect 75680 26438 75728 26502
rect 75792 26438 75850 26502
rect 75680 26390 75850 26438
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect 551331 10581 551453 10587
rect 551331 10464 551336 10469
rect 551448 10464 551453 10469
rect 551331 10459 551453 10464
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect 576153 9741 576275 9747
rect 576153 9624 576158 9629
rect 576270 9624 576275 9629
rect 576153 9619 576275 9624
rect -800 8636 480 8748
rect 69759 8651 69881 8657
rect 583520 8636 584800 8748
rect 69759 8534 69764 8539
rect 69876 8534 69881 8539
rect 69759 8529 69881 8534
rect 558423 7881 558545 7887
rect 558423 7764 558428 7769
rect 558540 7764 558545 7769
rect 558423 7759 558545 7764
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect 66359 7091 66481 7097
rect 66359 6974 66364 6979
rect 66476 6974 66481 6979
rect 66359 6969 66481 6974
rect 572607 6561 572729 6567
rect 572607 6444 572612 6449
rect 572724 6444 572729 6449
rect 572607 6439 572729 6444
rect -800 6272 480 6384
rect 565515 6311 565637 6317
rect 565515 6194 565520 6199
rect 565632 6194 565637 6199
rect 565515 6189 565637 6194
rect 569061 6291 569183 6297
rect 583520 6272 584800 6384
rect 569061 6174 569066 6179
rect 569178 6174 569183 6179
rect 569061 6169 569183 6174
rect 554877 6161 554999 6167
rect 554877 6044 554882 6049
rect 554994 6044 554999 6049
rect 554877 6039 554999 6044
rect 561969 6081 562091 6087
rect 561969 5964 561974 5969
rect 562086 5964 562091 5969
rect 561969 5959 562091 5964
rect 62869 5711 62991 5717
rect 62869 5594 62874 5599
rect 62986 5594 62991 5599
rect 62869 5589 62991 5594
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect 55239 4381 55361 4387
rect 55239 4264 55244 4269
rect 55356 4264 55361 4269
rect 55239 4259 55361 4264
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect 52329 3351 52451 3357
rect 52329 3234 52334 3239
rect 52446 3234 52451 3239
rect 52329 3229 52451 3234
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect 49529 2271 49651 2277
rect 49529 2154 49534 2159
rect 49646 2154 49651 2159
rect 49529 2149 49651 2154
rect 46409 1731 46531 1737
rect -800 1544 480 1656
rect 46409 1614 46414 1619
rect 46526 1614 46531 1619
rect 46409 1609 46531 1614
rect 583520 1544 584800 1656
<< via3 >>
rect 22590 695320 23050 695780
rect 23590 695310 24050 695770
rect 24590 695420 25050 695880
rect 25590 695420 26050 695880
rect 165595 699685 168093 699689
rect 165595 697195 165599 699685
rect 165599 697195 168089 699685
rect 168089 697195 168093 699685
rect 165595 697191 168093 697195
rect 218481 697631 220979 700129
rect 319171 698681 321669 701179
rect 26658 682328 26663 683627
rect 26663 682328 27687 683627
rect 27687 682328 27692 683627
rect 29711 682806 29716 683670
rect 29716 682806 30585 683670
rect 30585 682806 30590 683670
rect 31106 683151 31111 683644
rect 31111 683151 31609 683644
rect 31609 683151 31614 683644
rect 31106 683146 31614 683151
rect 29711 682801 30590 682806
rect 26658 682323 27692 682328
rect 22490 677810 24950 680270
rect 19000 634750 21460 637210
rect 14060 559600 16520 562060
rect 14400 549750 16860 552210
rect 40191 689345 42649 689349
rect 40191 686895 40195 689345
rect 40195 686895 42645 689345
rect 42645 686895 42649 689345
rect 40191 686891 42649 686895
rect 36783 295420 36895 295532
rect 29956 249971 30024 250039
rect 32588 206138 32652 206142
rect 32588 206082 32592 206138
rect 32592 206082 32648 206138
rect 32648 206082 32652 206138
rect 32588 206078 32652 206082
rect 24950 203217 26591 204858
rect 49575 204410 49645 204415
rect 49575 204351 49580 204410
rect 49580 204351 49640 204410
rect 49640 204351 49645 204410
rect 54111 211900 54175 211905
rect 54111 211840 54170 211900
rect 54170 211840 54175 211900
rect 54111 211835 54175 211840
rect 54510 209920 54574 209925
rect 54510 209860 54569 209920
rect 54569 209860 54574 209920
rect 54510 209855 54574 209860
rect 54945 207540 55009 207545
rect 54945 207480 55004 207540
rect 55004 207480 55009 207540
rect 54945 207475 55009 207480
rect 56525 205690 56595 205695
rect 56525 205631 56530 205690
rect 56530 205631 56590 205690
rect 56590 205631 56595 205690
rect 51752 202962 51816 203026
rect 53498 202998 53562 203002
rect 53498 202942 53502 202998
rect 53502 202942 53558 202998
rect 53558 202942 53562 202998
rect 53498 202938 53562 202942
rect 54838 202968 54902 202972
rect 54838 202912 54842 202968
rect 54842 202912 54898 202968
rect 54898 202912 54902 202968
rect 54838 202908 54902 202912
rect 55528 202948 55592 202952
rect 55528 202892 55532 202948
rect 55532 202892 55588 202948
rect 55588 202892 55592 202948
rect 55528 202888 55592 202892
rect 54227 202858 54291 202862
rect 54227 202802 54231 202858
rect 54231 202802 54287 202858
rect 54287 202802 54291 202858
rect 54227 202798 54291 202802
rect 44915 201070 45215 201075
rect 44915 200770 44920 201070
rect 44920 200770 45215 201070
rect 44915 200765 45215 200770
rect 24649 199640 25774 200765
rect 45015 200130 45315 200135
rect 45015 199830 45020 200130
rect 45020 199830 45315 200130
rect 45015 199825 45315 199830
rect 49184 199490 49254 199560
rect 45445 199110 45745 199115
rect 45445 198810 45450 199110
rect 45450 198810 45745 199110
rect 45445 198805 45745 198810
rect 24781 195324 27241 197784
rect 55765 196350 55865 196355
rect 55765 196250 55860 196350
rect 55860 196250 55865 196350
rect 55765 196245 55865 196250
rect 24930 188852 27390 191312
rect 24639 182507 27099 184967
rect 75728 26498 75792 26502
rect 75728 26442 75732 26498
rect 75732 26442 75788 26498
rect 75788 26442 75792 26498
rect 75728 26438 75792 26442
rect 551331 10576 551453 10581
rect 551331 10469 551336 10576
rect 551336 10469 551448 10576
rect 551448 10469 551453 10576
rect 576153 9736 576275 9741
rect 576153 9629 576158 9736
rect 576158 9629 576270 9736
rect 576270 9629 576275 9736
rect 69759 8646 69881 8651
rect 69759 8539 69764 8646
rect 69764 8539 69876 8646
rect 69876 8539 69881 8646
rect 558423 7876 558545 7881
rect 558423 7769 558428 7876
rect 558428 7769 558540 7876
rect 558540 7769 558545 7876
rect 66359 7086 66481 7091
rect 66359 6979 66364 7086
rect 66364 6979 66476 7086
rect 66476 6979 66481 7086
rect 572607 6556 572729 6561
rect 572607 6449 572612 6556
rect 572612 6449 572724 6556
rect 572724 6449 572729 6556
rect 565515 6306 565637 6311
rect 565515 6199 565520 6306
rect 565520 6199 565632 6306
rect 565632 6199 565637 6306
rect 569061 6286 569183 6291
rect 569061 6179 569066 6286
rect 569066 6179 569178 6286
rect 569178 6179 569183 6286
rect 554877 6156 554999 6161
rect 554877 6049 554882 6156
rect 554882 6049 554994 6156
rect 554994 6049 554999 6156
rect 561969 6076 562091 6081
rect 561969 5969 561974 6076
rect 561974 5969 562086 6076
rect 562086 5969 562091 6076
rect 62869 5706 62991 5711
rect 62869 5599 62874 5706
rect 62874 5599 62986 5706
rect 62986 5599 62991 5706
rect 55239 4376 55361 4381
rect 55239 4269 55244 4376
rect 55244 4269 55356 4376
rect 55356 4269 55361 4376
rect 52329 3346 52451 3351
rect 52329 3239 52334 3346
rect 52334 3239 52446 3346
rect 52446 3239 52451 3346
rect 49529 2266 49651 2271
rect 49529 2159 49534 2266
rect 49534 2159 49646 2266
rect 49646 2159 49651 2266
rect 46409 1726 46531 1731
rect 46409 1619 46414 1726
rect 46414 1619 46526 1726
rect 46526 1619 46531 1726
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 165594 699689 168094 702300
rect 165594 697191 165595 699689
rect 168093 697191 168094 699689
rect 218480 700129 220980 702300
rect 218480 697631 218481 700129
rect 220979 697631 220980 700129
rect 218480 697630 220980 697631
rect 319170 701179 321670 702300
rect 319170 698681 319171 701179
rect 321669 698681 321670 701179
rect 165594 697190 168094 697191
rect 319170 696530 321670 698681
rect 23049 695780 23051 695781
rect 23050 695320 23051 695780
rect 23049 695319 23051 695320
rect 20970 691430 42990 693890
rect 20970 684190 23430 691430
rect 40190 690040 42650 691430
rect 35930 689349 42910 690040
rect 35930 686891 40191 689349
rect 42649 686891 42910 689349
rect 35930 686320 42910 686891
rect 40190 684190 42650 686320
rect 20970 683670 42650 684190
rect 20970 683627 29711 683670
rect 20970 682323 26658 683627
rect 27692 682801 29711 683627
rect 30590 683644 42650 683670
rect 30590 683146 31106 683644
rect 31614 683146 42650 683644
rect 30590 682801 42650 683146
rect 27692 682323 42650 682801
rect 20970 681730 42650 682323
rect 22489 680270 22491 680271
rect 22489 677810 22490 680270
rect 22489 677809 22491 677810
rect 18999 637210 19001 637211
rect 18999 634750 19000 637210
rect 18999 634749 19001 634750
rect 14059 562060 16521 562061
rect 36140 562060 38600 681730
rect 40190 562060 42650 681730
rect 14059 559600 14060 562060
rect 16520 559600 44190 562060
rect 14059 559599 16521 559600
rect 14399 552210 16861 552211
rect 24506 552210 26966 559600
rect 36140 552210 38600 559600
rect 14399 549750 14400 552210
rect 16860 549750 38600 552210
rect 14399 549749 16861 549750
rect 24506 204858 26966 549750
rect 36829 295533 36889 297140
rect 36782 295532 36896 295533
rect 36782 295420 36783 295532
rect 36895 295420 36896 295532
rect 36782 295419 36896 295420
rect 24506 203217 24950 204858
rect 26591 203217 26966 204858
rect 24506 200765 26966 203217
rect 24506 199640 24649 200765
rect 25774 199640 26966 200765
rect 24506 197785 26966 199640
rect 29955 250039 30025 250040
rect 29955 249971 29956 250039
rect 30024 249971 30025 250039
rect 29955 199560 30025 249971
rect 36829 209382 36889 295419
rect 36829 209322 50973 209382
rect 32587 206142 32653 206143
rect 32587 206078 32588 206142
rect 32652 206140 32653 206142
rect 49580 206140 49640 206350
rect 32652 206080 49640 206140
rect 32652 206078 32653 206080
rect 32587 206077 32653 206078
rect 49580 204416 49640 206080
rect 49574 204415 49646 204416
rect 49574 204351 49575 204415
rect 49645 204351 49646 204415
rect 49574 204350 49646 204351
rect 50913 202301 50973 209322
rect 53510 207580 53570 213020
rect 54020 210237 54080 210740
rect 54020 210177 54298 210237
rect 54020 210077 54080 210177
rect 54238 208290 54298 210177
rect 54211 208230 54479 208290
rect 54238 208223 54298 208230
rect 53984 207580 54044 207688
rect 53510 207520 54044 207580
rect 53510 207488 53570 207520
rect 53984 204790 54044 207520
rect 54419 204750 54479 208230
rect 54640 207000 54700 208520
rect 54640 206940 54914 207000
rect 54854 204750 54914 206940
rect 55289 204750 55349 206470
rect 51751 203026 51817 203027
rect 51751 202962 51752 203026
rect 51816 202962 51817 203026
rect 51751 202961 51817 202962
rect 53497 203002 53563 203003
rect 51754 202301 51814 202961
rect 53497 202938 53498 203002
rect 53562 203000 53563 203002
rect 53794 203000 53854 203130
rect 53562 202940 53854 203000
rect 53562 202938 53563 202940
rect 53497 202937 53563 202938
rect 54229 202863 54289 203120
rect 54664 202970 54724 203110
rect 54837 202972 54903 202973
rect 54837 202970 54838 202972
rect 54664 202910 54838 202970
rect 54837 202908 54838 202910
rect 54902 202908 54903 202972
rect 54837 202907 54903 202908
rect 55099 202950 55159 203110
rect 55527 202952 55593 202953
rect 55527 202950 55528 202952
rect 55099 202890 55528 202950
rect 55527 202888 55528 202890
rect 55592 202950 55593 202952
rect 55592 202890 55600 202950
rect 55592 202888 55593 202890
rect 55527 202887 55593 202888
rect 54226 202862 54292 202863
rect 54226 202798 54227 202862
rect 54291 202798 54292 202862
rect 54226 202797 54292 202798
rect 50913 202241 51814 202301
rect 44914 201075 45216 201076
rect 44914 200765 44915 201075
rect 45215 200765 45216 201075
rect 44914 200764 45216 200765
rect 45014 200135 45316 200136
rect 45014 199825 45015 200135
rect 45315 199825 45316 200135
rect 45014 199824 45316 199825
rect 49183 199560 49255 199561
rect 29955 199490 49184 199560
rect 49254 199490 49255 199560
rect 49183 199489 49255 199490
rect 45444 199115 45746 199116
rect 45444 198805 45445 199115
rect 45745 198805 45746 199115
rect 45444 198804 45746 198805
rect 24506 197784 27242 197785
rect 24506 195324 24781 197784
rect 27241 195324 27242 197784
rect 24506 195323 27242 195324
rect 24506 191313 26966 195323
rect 24506 191312 27391 191313
rect 24506 188852 24930 191312
rect 27390 188852 27391 191312
rect 24506 188851 27391 188852
rect 24506 184968 26966 188851
rect 24506 184967 27100 184968
rect 24506 182507 24639 184967
rect 27099 182507 27100 184967
rect 24506 182506 27100 182507
rect 24506 181365 26966 182506
rect 46414 13050 46526 13066
rect 53050 13050 53110 198800
rect 45470 12990 53110 13050
rect 46414 1732 46526 12990
rect 49534 11770 49646 11956
rect 53390 11770 53450 198800
rect 48760 11710 53450 11770
rect 49534 2272 49646 11710
rect 52334 6940 52446 7926
rect 53730 6940 53790 198800
rect 54070 11260 54130 198800
rect 54410 15140 54470 198800
rect 54750 19490 54810 198800
rect 55090 25220 55150 198800
rect 55430 26500 55490 198800
rect 55764 196355 55866 196356
rect 55764 196245 55765 196355
rect 55865 196245 55866 196355
rect 55764 196244 55866 196245
rect 75727 26502 75793 26503
rect 75727 26500 75728 26502
rect 55430 26440 75728 26500
rect 75727 26438 75728 26440
rect 75792 26438 75793 26502
rect 75727 26437 75793 26438
rect 69764 25220 69876 25276
rect 55090 25160 70080 25220
rect 66364 19490 66476 19546
rect 54750 19430 67040 19490
rect 62874 15140 62986 15746
rect 54410 15080 63110 15140
rect 55244 11260 55356 11286
rect 54070 11200 58680 11260
rect 51770 6880 53790 6940
rect 52334 3352 52446 6880
rect 53730 6770 53790 6880
rect 55244 4382 55356 11200
rect 62874 5712 62986 15080
rect 66364 7092 66476 19430
rect 69764 8652 69876 25160
rect 69758 8651 69882 8652
rect 69758 8539 69759 8651
rect 69881 8539 69882 8651
rect 69758 8538 69882 8539
rect 66358 7091 66482 7092
rect 66358 6979 66359 7091
rect 66481 6979 66482 7091
rect 66358 6978 66482 6979
rect 62868 5711 62992 5712
rect 62868 5599 62869 5711
rect 62991 5599 62992 5711
rect 62868 5598 62992 5599
rect 55238 4381 55362 4382
rect 55238 4269 55239 4381
rect 55361 4269 55362 4381
rect 55238 4268 55362 4269
rect 52328 3351 52452 3352
rect 52328 3239 52329 3351
rect 52451 3239 52452 3351
rect 52328 3238 52452 3239
rect 49528 2271 49652 2272
rect 49528 2159 49529 2271
rect 49651 2159 49652 2271
rect 49528 2158 49652 2159
rect 46408 1731 46532 1732
rect 46408 1619 46409 1731
rect 46531 1619 46532 1731
rect 46408 1618 46532 1619
<< via4 >>
rect 24589 695880 25051 695881
rect 22589 695780 23049 695781
rect 22589 695320 22590 695780
rect 22590 695320 23049 695780
rect 22589 695319 23049 695320
rect 23589 695770 24051 695771
rect 23589 695310 23590 695770
rect 23590 695310 24050 695770
rect 24050 695310 24051 695770
rect 24589 695420 24590 695880
rect 24590 695420 25050 695880
rect 25050 695420 25051 695880
rect 24589 695419 25051 695420
rect 25589 695880 26051 695881
rect 25589 695420 25590 695880
rect 25590 695420 26050 695880
rect 26050 695420 26051 695880
rect 25589 695419 26051 695420
rect 23589 695309 24051 695310
rect 22491 680270 24951 680271
rect 22491 677810 24950 680270
rect 24950 677810 24951 680270
rect 22491 677809 24951 677810
rect 19001 637210 21461 637211
rect 19001 634750 21460 637210
rect 21460 634750 21461 637210
rect 19001 634749 21461 634750
rect 53380 213020 53700 213340
rect 53983 211905 54303 212030
rect 53983 211835 54111 211905
rect 54111 211835 54175 211905
rect 54175 211835 54303 211905
rect 53983 211710 54303 211835
rect 53890 210740 54210 211060
rect 54382 209925 54702 210050
rect 54382 209855 54510 209925
rect 54510 209855 54574 209925
rect 54574 209855 54702 209925
rect 54382 209730 54702 209855
rect 54510 208520 54830 208840
rect 54817 207545 55137 207670
rect 54817 207475 54945 207545
rect 54945 207475 55009 207545
rect 55009 207475 55137 207545
rect 54817 207350 55137 207475
rect 55159 206470 55479 206790
rect 56400 205695 56720 205823
rect 56400 205631 56525 205695
rect 56525 205631 56595 205695
rect 56595 205631 56720 205695
rect 56400 205503 56720 205631
rect 551232 10581 551552 10685
rect 551232 10469 551331 10581
rect 551331 10469 551453 10581
rect 551453 10469 551552 10581
rect 551232 10365 551552 10469
rect 576054 9741 576374 9845
rect 576054 9629 576153 9741
rect 576153 9629 576275 9741
rect 576275 9629 576374 9741
rect 576054 9525 576374 9629
rect 558324 7881 558644 7985
rect 558324 7769 558423 7881
rect 558423 7769 558545 7881
rect 558545 7769 558644 7881
rect 558324 7665 558644 7769
rect 572508 6561 572828 6665
rect 572508 6449 572607 6561
rect 572607 6449 572729 6561
rect 572729 6449 572828 6561
rect 565416 6311 565736 6415
rect 554778 6161 555098 6265
rect 565416 6199 565515 6311
rect 565515 6199 565637 6311
rect 565637 6199 565736 6311
rect 554778 6049 554877 6161
rect 554877 6049 554999 6161
rect 554999 6049 555098 6161
rect 554778 5945 555098 6049
rect 561870 6081 562190 6185
rect 565416 6095 565736 6199
rect 568962 6291 569282 6395
rect 572508 6345 572828 6449
rect 568962 6179 569061 6291
rect 569061 6179 569183 6291
rect 569183 6179 569282 6291
rect 561870 5969 561969 6081
rect 561969 5969 562091 6081
rect 562091 5969 562190 6081
rect 568962 6075 569282 6179
rect 561870 5865 562190 5969
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 16200 695881 52140 697010
rect 16200 695781 24589 695881
rect 16200 695319 22589 695781
rect 23049 695771 24589 695781
rect 23049 695319 23589 695771
rect 16200 695309 23589 695319
rect 24051 695419 24589 695771
rect 25051 695419 25589 695881
rect 26051 695419 52140 695881
rect 24051 695309 52140 695419
rect 16200 694550 52140 695309
rect 16200 680270 18660 694550
rect 22467 680271 24975 680295
rect 22467 680270 22491 680271
rect 16200 677830 22491 680270
rect 16300 677810 22491 677830
rect 22467 677809 22491 677810
rect 24951 680270 24975 680271
rect 49680 680270 52140 694550
rect 24951 677810 52140 680270
rect 24951 677809 25340 677810
rect 22467 677785 25340 677809
rect 18977 637211 21485 637235
rect 18977 634749 19001 637211
rect 21461 637210 21485 637211
rect 22880 637210 25340 677785
rect 26710 637210 29170 677810
rect 21461 634750 29170 637210
rect 21461 634749 21485 634750
rect 18977 634725 21485 634749
rect 336440 234570 336760 235580
rect 336400 234250 576374 234570
rect 53356 213340 53724 213364
rect 336440 213340 336760 234250
rect 53356 213020 53380 213340
rect 53700 213020 336760 213340
rect 338550 229440 338870 230130
rect 572508 229440 572828 231090
rect 338550 229120 572828 229440
rect 53356 212996 53724 213020
rect 53959 212030 54327 212054
rect 338550 212030 338870 229120
rect 53959 211710 53983 212030
rect 54303 211710 338870 212030
rect 340730 226010 341050 226430
rect 340730 225690 569282 226010
rect 53959 211686 54327 211710
rect 53866 211060 54234 211084
rect 340730 211060 341050 225690
rect 342450 223150 342770 223950
rect 342380 222830 565736 223150
rect 53866 210740 53890 211060
rect 54210 210740 341050 211060
rect 53866 210716 54234 210740
rect 54358 210050 54726 210074
rect 342450 210050 342770 222830
rect 344410 220290 344730 220460
rect 344380 219970 562190 220290
rect 54358 209730 54382 210050
rect 54702 209730 342770 210050
rect 54358 209706 54726 209730
rect 54486 208840 54854 208864
rect 344410 208840 344730 219970
rect 54486 208520 54510 208840
rect 54830 208520 344730 208840
rect 346240 215530 346560 215810
rect 346240 215210 558644 215530
rect 54486 208496 54854 208520
rect 54793 207670 55161 207694
rect 346240 207670 346560 215210
rect 554778 211080 555098 212500
rect 354950 210760 555098 211080
rect 54793 207350 54817 207670
rect 55137 207350 346560 207670
rect 54793 207326 55161 207350
rect 55135 206790 55503 206814
rect 355080 206790 355400 210760
rect 356420 208920 551552 209240
rect 55135 206470 55159 206790
rect 55479 206470 355400 206790
rect 55135 206446 55503 206470
rect 56400 206050 56720 206060
rect 356460 206050 356780 208920
rect 56400 206020 356780 206050
rect 56330 205823 356780 206020
rect 56330 205503 56400 205823
rect 56720 205730 356780 205823
rect 56720 205503 56940 205730
rect 56330 205460 56940 205503
rect 551232 10709 551552 208920
rect 551208 10685 551576 10709
rect 551208 10365 551232 10685
rect 551552 10365 551576 10685
rect 551208 10341 551576 10365
rect 554778 6289 555098 210760
rect 558324 8009 558644 215210
rect 558300 7985 558668 8009
rect 558300 7665 558324 7985
rect 558644 7665 558668 7985
rect 558300 7641 558668 7665
rect 554754 6265 555122 6289
rect 554754 5945 554778 6265
rect 555098 5945 555122 6265
rect 561870 6209 562190 219970
rect 565416 6439 565736 222830
rect 565392 6415 565760 6439
rect 568962 6419 569282 225690
rect 572508 6689 572828 229120
rect 576054 226910 576374 234250
rect 573940 226590 576374 226910
rect 576054 9869 576374 226590
rect 576030 9845 576398 9869
rect 576030 9525 576054 9845
rect 576374 9525 576398 9845
rect 576030 9501 576398 9525
rect 572484 6665 572852 6689
rect 554754 5921 555122 5945
rect 561846 6185 562214 6209
rect 561846 5865 561870 6185
rect 562190 5865 562214 6185
rect 565392 6095 565416 6415
rect 565736 6095 565760 6415
rect 565392 6071 565760 6095
rect 568938 6395 569306 6419
rect 568938 6075 568962 6395
rect 569282 6075 569306 6395
rect 572484 6345 572508 6665
rect 572828 6345 572852 6665
rect 572484 6321 572852 6345
rect 568938 6051 569306 6075
rect 561846 5841 562214 5865
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use 8bit_sens  8bit_sens_0
timestamp 1661898952
transform 1 0 52880 0 1 199490
box -110 -750 2810 3340
use adc  adc_0
timestamp 1662015318
transform 1 0 52980 0 1 205530
box 450 -2480 2630 -665
use bias_cell  bias_cell_0
timestamp 1661984010
transform 1 0 24660 0 1 691160
box 790 -2240 11230 -60
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
