magic
tech sky130B
magscale 1 2
timestamp 1662180122
<< metal2 >>
rect 311 4155 320 4225
rect 390 4155 399 4225
rect 320 3485 390 4155
rect 450 3995 520 4250
rect 441 3925 450 3995
rect 520 3925 529 3995
rect 450 3500 520 3925
rect 680 3785 750 3794
rect 680 3495 750 3715
rect 1564 3507 1604 4370
rect 1999 3495 2039 4340
rect 2434 3527 2474 4370
rect 2869 3525 2909 4360
<< via2 >>
rect 320 4155 390 4225
rect 450 3925 520 3995
rect 680 3715 750 3785
<< metal3 >>
rect 60 4225 3560 4290
rect 60 4155 320 4225
rect 390 4155 3560 4225
rect 60 4110 3560 4155
rect 50 3995 3550 4050
rect 50 3925 450 3995
rect 520 3925 3560 3995
rect 50 3870 3550 3925
rect 50 3785 3550 3810
rect 50 3715 680 3785
rect 750 3715 3560 3785
rect 50 3630 3550 3715
<< metal4 >>
rect 1464 3502 1524 4360
rect 1899 3501 1959 4370
rect 2334 3510 2394 4380
rect 2769 3510 2829 4360
use pixel  pixel_0
timestamp 1662180122
transform 1 0 460 0 1 3000
box -470 -3000 3090 570
<< labels >>
rlabel metal2 2889 3739 2889 3739 1 GRAYx0x
port 1 n
rlabel metal4 2796 3759 2796 3759 1 GRAYx1x
port 2 n
rlabel metal2 2460 3780 2460 3780 1 GRAYx2x
port 3 n
rlabel metal4 2360 3760 2360 3760 1 GRAYx3x
port 4 n
rlabel metal2 2020 3740 2020 3740 1 GRAYx4x
port 5 n
rlabel metal4 1930 3740 1930 3740 1 GRAYx5x
port 6 n
rlabel metal2 1580 3760 1580 3760 1 GRAYx6x
port 7 n
rlabel metal4 1490 3760 1490 3760 1 GRAYx7x
port 8 n
<< end >>
