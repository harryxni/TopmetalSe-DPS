magic
tech sky130B
magscale 1 2
timestamp 1607692587
<< nwell >>
rect 0 370 1880 640
rect 0 298 474 370
rect 792 368 1880 370
rect 792 298 1020 368
rect 1334 320 1880 368
rect 1334 310 1572 320
rect 1372 296 1572 310
<< pwell >>
rect 6 30 90 64
rect 174 30 258 64
rect 334 30 418 64
rect 604 30 688 64
rect 788 30 872 64
rect 1000 30 1084 64
rect 1168 30 1252 64
rect 1404 30 1488 64
rect 1572 30 1656 64
rect 1740 30 1824 64
<< nmos >>
rect 128 134 158 222
rect 350 130 380 222
rect 634 134 664 302
rect 896 128 926 220
rect 1164 132 1194 300
rect 1442 130 1472 222
rect 1652 118 1682 210
rect 1754 118 1784 210
<< pmos >>
rect 128 346 158 490
rect 350 346 380 490
rect 634 408 664 492
rect 896 344 926 488
rect 1164 406 1194 490
rect 1442 346 1472 490
rect 1652 366 1682 510
rect 1754 366 1784 510
<< ndiff >>
rect 576 284 634 302
rect 576 250 588 284
rect 622 250 634 284
rect 70 204 128 222
rect 70 170 82 204
rect 116 170 128 204
rect 70 134 128 170
rect 158 204 216 222
rect 158 170 170 204
rect 204 170 216 204
rect 158 134 216 170
rect 290 204 350 222
rect 290 170 304 204
rect 338 170 350 204
rect 290 130 350 170
rect 380 204 438 222
rect 380 170 392 204
rect 426 170 438 204
rect 576 216 634 250
rect 380 130 438 170
rect 576 182 588 216
rect 622 182 634 216
rect 576 134 634 182
rect 664 284 722 302
rect 664 250 676 284
rect 710 250 722 284
rect 664 216 722 250
rect 1106 282 1164 300
rect 1106 248 1118 282
rect 1152 248 1164 282
rect 664 182 676 216
rect 710 182 722 216
rect 664 134 722 182
rect 838 202 896 220
rect 838 168 850 202
rect 884 168 896 202
rect 838 128 896 168
rect 926 202 984 220
rect 926 168 938 202
rect 972 168 984 202
rect 1106 214 1164 248
rect 926 128 984 168
rect 1106 180 1118 214
rect 1152 180 1164 214
rect 1106 132 1164 180
rect 1194 282 1252 300
rect 1194 248 1206 282
rect 1240 248 1252 282
rect 1194 214 1252 248
rect 1194 180 1206 214
rect 1240 180 1252 214
rect 1194 132 1252 180
rect 1384 204 1442 222
rect 1384 170 1396 204
rect 1430 170 1442 204
rect 1384 130 1442 170
rect 1472 204 1530 222
rect 1472 170 1484 204
rect 1518 170 1530 204
rect 1472 130 1530 170
rect 1590 176 1652 210
rect 1590 142 1602 176
rect 1636 142 1652 176
rect 1590 118 1652 142
rect 1682 166 1754 210
rect 1682 132 1706 166
rect 1740 132 1754 166
rect 1682 118 1754 132
rect 1784 176 1842 210
rect 1784 142 1800 176
rect 1834 142 1842 176
rect 1784 118 1842 142
<< pdiff >>
rect 70 482 128 490
rect 70 448 82 482
rect 116 448 128 482
rect 70 414 128 448
rect 70 380 82 414
rect 116 380 128 414
rect 70 346 128 380
rect 158 456 216 490
rect 158 422 170 456
rect 204 422 216 456
rect 158 388 216 422
rect 158 354 170 388
rect 204 354 216 388
rect 158 346 216 354
rect 292 482 350 490
rect 292 448 304 482
rect 338 448 350 482
rect 292 414 350 448
rect 292 380 304 414
rect 338 380 350 414
rect 292 346 350 380
rect 380 456 438 490
rect 380 422 392 456
rect 426 422 438 456
rect 576 466 634 492
rect 380 388 438 422
rect 576 432 588 466
rect 622 432 634 466
rect 576 408 634 432
rect 664 464 722 492
rect 664 430 676 464
rect 710 430 722 464
rect 664 408 722 430
rect 838 480 896 488
rect 838 446 850 480
rect 884 446 896 480
rect 838 412 896 446
rect 380 354 392 388
rect 426 354 438 388
rect 380 346 438 354
rect 838 378 850 412
rect 884 378 896 412
rect 838 344 896 378
rect 926 454 984 488
rect 926 420 938 454
rect 972 420 984 454
rect 926 386 984 420
rect 1106 464 1164 490
rect 1106 430 1118 464
rect 1152 430 1164 464
rect 1106 406 1164 430
rect 1194 462 1252 490
rect 1194 428 1206 462
rect 1240 428 1252 462
rect 1590 502 1652 510
rect 1384 482 1442 490
rect 1384 448 1396 482
rect 1430 448 1442 482
rect 1194 406 1252 428
rect 1384 414 1442 448
rect 926 352 938 386
rect 972 352 984 386
rect 1384 380 1396 414
rect 1430 380 1442 414
rect 926 344 984 352
rect 1384 346 1442 380
rect 1472 456 1530 490
rect 1472 422 1484 456
rect 1518 422 1530 456
rect 1472 388 1530 422
rect 1472 354 1484 388
rect 1518 354 1530 388
rect 1590 468 1602 502
rect 1636 468 1652 502
rect 1590 434 1652 468
rect 1590 400 1602 434
rect 1636 400 1652 434
rect 1590 366 1652 400
rect 1682 502 1754 510
rect 1682 468 1704 502
rect 1738 468 1754 502
rect 1682 366 1754 468
rect 1784 502 1844 510
rect 1784 468 1798 502
rect 1832 468 1844 502
rect 1784 434 1844 468
rect 1784 400 1798 434
rect 1832 400 1844 434
rect 1784 366 1842 400
rect 1472 346 1530 354
<< ndiffc >>
rect 588 250 622 284
rect 82 170 116 204
rect 170 170 204 204
rect 304 170 338 204
rect 392 170 426 204
rect 588 182 622 216
rect 676 250 710 284
rect 1118 248 1152 282
rect 676 182 710 216
rect 850 168 884 202
rect 938 168 972 202
rect 1118 180 1152 214
rect 1206 248 1240 282
rect 1206 180 1240 214
rect 1396 170 1430 204
rect 1484 170 1518 204
rect 1602 142 1636 176
rect 1706 132 1740 166
rect 1800 142 1834 176
<< pdiffc >>
rect 82 448 116 482
rect 82 380 116 414
rect 170 422 204 456
rect 170 354 204 388
rect 304 448 338 482
rect 304 380 338 414
rect 392 422 426 456
rect 588 432 622 466
rect 676 430 710 464
rect 850 446 884 480
rect 392 354 426 388
rect 850 378 884 412
rect 938 420 972 454
rect 1118 430 1152 464
rect 1206 428 1240 462
rect 1396 448 1430 482
rect 938 352 972 386
rect 1396 380 1430 414
rect 1484 422 1518 456
rect 1484 354 1518 388
rect 1602 468 1636 502
rect 1602 400 1636 434
rect 1704 468 1738 502
rect 1798 468 1832 502
rect 1798 400 1832 434
<< psubdiff >>
rect 6 30 32 64
rect 66 30 90 64
rect 174 30 200 64
rect 234 30 258 64
rect 334 30 360 64
rect 394 30 418 64
rect 604 30 630 64
rect 664 30 688 64
rect 788 30 814 64
rect 848 30 872 64
rect 1000 30 1026 64
rect 1060 30 1084 64
rect 1168 30 1194 64
rect 1228 30 1252 64
rect 1404 30 1430 64
rect 1464 30 1488 64
rect 1572 30 1598 64
rect 1632 30 1656 64
rect 1740 30 1766 64
rect 1800 30 1824 64
<< nsubdiff >>
rect 86 602 172 604
rect 86 568 112 602
rect 146 568 172 602
rect 86 566 172 568
rect 250 602 336 604
rect 250 568 276 602
rect 310 568 336 602
rect 250 566 336 568
rect 540 602 626 604
rect 540 568 566 602
rect 600 568 626 602
rect 540 566 626 568
rect 696 602 782 604
rect 696 568 722 602
rect 756 568 782 602
rect 696 566 782 568
rect 884 602 970 604
rect 884 568 910 602
rect 944 568 970 602
rect 884 566 970 568
rect 1100 602 1186 604
rect 1100 568 1126 602
rect 1160 568 1186 602
rect 1100 566 1186 568
rect 1340 602 1426 604
rect 1340 568 1366 602
rect 1400 568 1426 602
rect 1340 566 1426 568
rect 1512 602 1598 604
rect 1512 568 1538 602
rect 1572 568 1598 602
rect 1512 566 1598 568
rect 1684 602 1770 604
rect 1684 568 1710 602
rect 1744 568 1770 602
rect 1684 566 1770 568
<< psubdiffcont >>
rect 32 30 66 64
rect 200 30 234 64
rect 360 30 394 64
rect 630 30 664 64
rect 814 30 848 64
rect 1026 30 1060 64
rect 1194 30 1228 64
rect 1430 30 1464 64
rect 1598 30 1632 64
rect 1766 30 1800 64
<< nsubdiffcont >>
rect 112 568 146 602
rect 276 568 310 602
rect 566 568 600 602
rect 722 568 756 602
rect 910 568 944 602
rect 1126 568 1160 602
rect 1366 568 1400 602
rect 1538 568 1572 602
rect 1710 568 1744 602
<< poly >>
rect 128 490 158 516
rect 350 490 380 516
rect 478 514 664 544
rect 478 494 532 514
rect 478 460 488 494
rect 522 460 532 494
rect 634 492 664 514
rect 478 444 532 460
rect 896 488 926 514
rect 1164 512 1344 542
rect 1164 490 1194 512
rect 634 380 664 408
rect 128 306 158 346
rect 350 306 380 346
rect 1290 482 1344 512
rect 1442 490 1472 516
rect 1652 510 1682 536
rect 1754 510 1784 536
rect 1290 448 1300 482
rect 1334 448 1344 482
rect 1290 432 1344 448
rect 1164 378 1194 406
rect 70 302 158 306
rect 292 302 380 306
rect 634 302 664 328
rect 896 304 926 344
rect 64 296 158 302
rect 64 262 82 296
rect 116 262 158 296
rect 64 254 158 262
rect 286 296 380 302
rect 286 262 304 296
rect 338 262 380 296
rect 286 254 380 262
rect 70 252 158 254
rect 292 252 380 254
rect 128 222 158 252
rect 350 222 380 252
rect 128 108 158 134
rect 480 184 534 200
rect 480 150 490 184
rect 524 150 534 184
rect 350 104 380 130
rect 480 118 534 150
rect 838 300 926 304
rect 1164 300 1194 326
rect 1442 306 1472 346
rect 1652 334 1682 366
rect 1754 336 1784 366
rect 1384 302 1472 306
rect 832 294 926 300
rect 832 260 850 294
rect 884 260 926 294
rect 832 252 926 260
rect 838 250 926 252
rect 896 220 926 250
rect 634 118 664 134
rect 1024 176 1078 192
rect 1024 142 1034 176
rect 1068 142 1078 176
rect 480 88 664 118
rect 896 102 926 128
rect 1024 116 1078 142
rect 1378 296 1472 302
rect 1378 262 1396 296
rect 1430 262 1472 296
rect 1620 318 1682 334
rect 1748 328 1784 336
rect 1620 284 1636 318
rect 1670 284 1684 318
rect 1726 310 1784 328
rect 1620 268 1682 284
rect 1378 254 1472 262
rect 1384 252 1472 254
rect 1442 222 1472 252
rect 1164 116 1194 132
rect 1652 210 1682 268
rect 1726 276 1736 310
rect 1770 276 1784 310
rect 1726 260 1784 276
rect 1748 248 1784 260
rect 1754 210 1784 248
rect 1024 86 1194 116
rect 1442 104 1472 130
rect 1652 92 1682 118
rect 1754 92 1784 118
<< polycont >>
rect 488 460 522 494
rect 1300 448 1334 482
rect 82 262 116 296
rect 304 262 338 296
rect 490 150 524 184
rect 850 260 884 294
rect 1034 142 1068 176
rect 1396 262 1430 296
rect 1636 284 1670 318
rect 1736 276 1770 310
<< locali >>
rect 0 602 1864 604
rect 0 568 112 602
rect 146 568 276 602
rect 310 568 566 602
rect 600 568 722 602
rect 756 568 910 602
rect 944 568 1126 602
rect 1160 568 1366 602
rect 1400 568 1538 602
rect 1572 568 1710 602
rect 1744 568 1864 602
rect 0 566 1864 568
rect 82 482 116 566
rect 82 414 116 448
rect 82 346 116 380
rect 170 456 204 490
rect 170 388 204 422
rect 170 312 204 354
rect 304 482 338 566
rect 488 494 522 510
rect 304 414 338 448
rect 304 346 338 380
rect 392 456 426 490
rect 488 444 522 459
rect 588 466 622 492
rect 392 388 426 422
rect 588 386 622 432
rect 392 314 426 354
rect 478 326 622 386
rect 478 314 528 326
rect 170 298 230 312
rect 0 262 82 296
rect 116 262 132 296
rect 170 264 182 298
rect 216 264 230 298
rect 170 252 230 264
rect 286 262 304 296
rect 338 262 354 296
rect 392 254 528 314
rect 588 284 622 326
rect 82 204 116 222
rect 82 64 116 170
rect 170 204 204 252
rect 170 150 204 170
rect 304 204 338 222
rect 304 64 338 170
rect 392 204 426 254
rect 588 216 622 250
rect 392 150 426 170
rect 474 150 490 184
rect 524 150 540 184
rect 588 166 622 182
rect 676 464 710 492
rect 676 380 710 430
rect 850 480 884 566
rect 850 412 884 446
rect 676 326 816 380
rect 850 344 884 378
rect 938 454 972 488
rect 938 386 972 420
rect 1118 464 1152 490
rect 1118 382 1152 430
rect 676 284 710 326
rect 782 308 816 326
rect 938 312 972 352
rect 1018 324 1152 382
rect 1018 312 1074 324
rect 782 304 824 308
rect 782 294 892 304
rect 782 260 850 294
rect 884 260 900 294
rect 782 254 892 260
rect 938 254 1074 312
rect 1118 282 1152 324
rect 676 216 710 250
rect 676 166 710 182
rect 850 202 884 220
rect 474 148 540 150
rect 850 64 884 168
rect 938 202 972 254
rect 1118 214 1152 248
rect 938 148 972 168
rect 1018 142 1034 176
rect 1068 142 1084 176
rect 1118 164 1152 180
rect 1206 462 1240 490
rect 1300 482 1334 500
rect 1300 432 1334 448
rect 1396 482 1430 566
rect 1596 502 1640 518
rect 1206 376 1240 428
rect 1396 414 1430 448
rect 1206 326 1314 376
rect 1396 346 1430 380
rect 1484 456 1518 490
rect 1484 388 1518 422
rect 1596 468 1602 502
rect 1636 468 1640 502
rect 1596 434 1640 468
rect 1698 502 1744 566
rect 1698 468 1704 502
rect 1738 468 1744 502
rect 1698 444 1744 468
rect 1798 510 1834 518
rect 1798 502 1856 510
rect 1832 468 1856 502
rect 1596 400 1602 434
rect 1636 402 1640 434
rect 1798 434 1856 468
rect 1636 400 1764 402
rect 1596 368 1764 400
rect 1206 282 1240 326
rect 1206 214 1240 248
rect 1206 164 1240 180
rect 1276 304 1314 326
rect 1484 312 1518 354
rect 1726 328 1764 368
rect 1832 400 1856 434
rect 1798 362 1856 400
rect 1806 328 1856 362
rect 1372 304 1438 306
rect 1276 296 1438 304
rect 1484 298 1552 312
rect 1276 262 1396 296
rect 1430 262 1446 296
rect 1484 264 1502 298
rect 1536 264 1552 298
rect 1618 284 1636 318
rect 1670 284 1686 318
rect 1726 310 1770 328
rect 1726 276 1736 310
rect 1726 270 1770 276
rect 1276 256 1438 262
rect 1276 202 1314 256
rect 1484 252 1552 264
rect 1724 260 1770 270
rect 1396 204 1430 222
rect 1276 188 1332 202
rect 1276 154 1292 188
rect 1326 154 1332 188
rect 1276 140 1332 154
rect 1396 64 1430 170
rect 1484 204 1518 252
rect 1724 250 1760 260
rect 1484 150 1518 170
rect 1594 216 1760 250
rect 1594 176 1638 216
rect 1822 196 1856 328
rect 1594 142 1602 176
rect 1636 142 1638 176
rect 1594 124 1638 142
rect 1700 166 1744 182
rect 1700 132 1706 166
rect 1740 132 1744 166
rect 1700 64 1744 132
rect 1796 176 1856 196
rect 1796 142 1800 176
rect 1834 142 1856 176
rect 1796 124 1856 142
rect 0 30 32 64
rect 66 30 200 64
rect 234 30 360 64
rect 394 30 630 64
rect 664 30 814 64
rect 848 30 1026 64
rect 1060 30 1194 64
rect 1228 30 1430 64
rect 1464 30 1598 64
rect 1632 30 1766 64
rect 1800 30 1870 64
<< viali >>
rect 112 568 146 602
rect 276 568 310 602
rect 566 568 600 602
rect 722 568 756 602
rect 910 568 944 602
rect 1126 568 1160 602
rect 1366 568 1400 602
rect 1538 568 1572 602
rect 1710 568 1744 602
rect 488 460 522 493
rect 488 459 522 460
rect 82 262 116 296
rect 182 264 216 298
rect 304 262 338 296
rect 490 150 524 184
rect 1034 142 1068 176
rect 1300 448 1334 482
rect 1502 264 1536 298
rect 1636 284 1670 318
rect 1292 154 1326 188
rect 32 30 66 64
rect 200 30 234 64
rect 360 30 394 64
rect 630 30 664 64
rect 814 30 848 64
rect 1026 30 1060 64
rect 1194 30 1228 64
rect 1430 30 1464 64
rect 1598 30 1632 64
rect 1766 30 1800 64
<< metal1 >>
rect 0 602 1864 640
rect 0 568 112 602
rect 146 568 276 602
rect 310 568 566 602
rect 600 568 722 602
rect 756 568 910 602
rect 944 568 1126 602
rect 1160 568 1366 602
rect 1400 568 1538 602
rect 1572 568 1710 602
rect 1744 568 1864 602
rect 0 544 1864 568
rect 474 502 538 508
rect 70 436 314 500
rect 474 450 480 502
rect 532 450 538 502
rect 1290 498 1346 500
rect 474 444 538 450
rect 1288 482 1346 498
rect 1288 448 1300 482
rect 1334 448 1346 482
rect 70 296 128 436
rect 264 414 314 436
rect 1288 432 1346 448
rect 1286 414 1344 432
rect 264 364 1344 414
rect 1624 318 1686 330
rect 70 262 82 296
rect 116 262 128 296
rect 70 254 128 262
rect 72 196 128 254
rect 166 310 236 318
rect 166 258 176 310
rect 228 258 236 310
rect 166 248 236 258
rect 292 298 1552 308
rect 292 296 1502 298
rect 292 262 304 296
rect 338 264 1502 296
rect 1536 264 1552 298
rect 1624 284 1636 318
rect 1670 284 1686 318
rect 1624 274 1686 284
rect 338 262 1552 264
rect 292 252 1552 262
rect 1630 200 1684 274
rect 72 184 542 196
rect 72 150 490 184
rect 524 150 542 184
rect 72 138 542 150
rect 1016 185 1082 192
rect 1016 133 1023 185
rect 1075 133 1082 185
rect 1280 188 1684 200
rect 1280 154 1292 188
rect 1326 154 1684 188
rect 1280 146 1684 154
rect 1280 142 1344 146
rect 1282 140 1344 142
rect 1016 126 1082 133
rect 0 64 1870 96
rect 0 30 32 64
rect 66 30 200 64
rect 234 30 360 64
rect 394 30 630 64
rect 664 30 814 64
rect 848 30 1026 64
rect 1060 30 1194 64
rect 1228 30 1430 64
rect 1464 30 1598 64
rect 1632 30 1766 64
rect 1800 30 1870 64
rect 0 0 1870 30
<< via1 >>
rect 480 493 532 502
rect 480 459 488 493
rect 488 459 522 493
rect 522 459 532 493
rect 480 450 532 459
rect 176 298 228 310
rect 176 264 182 298
rect 182 264 216 298
rect 216 264 228 298
rect 176 258 228 264
rect 1023 176 1075 185
rect 1023 142 1034 176
rect 1034 142 1068 176
rect 1068 142 1075 176
rect 1023 133 1075 142
<< metal2 >>
rect 474 450 480 502
rect 532 450 538 502
rect 170 318 236 332
rect 166 314 236 318
rect 474 314 538 450
rect 166 310 1080 314
rect 166 258 176 310
rect 228 258 1080 310
rect 166 256 1080 258
rect 166 248 236 256
rect 1014 186 1080 256
rect 1014 185 1082 186
rect 1014 174 1023 185
rect 1016 133 1023 174
rect 1075 133 1082 185
rect 1016 126 1082 133
<< labels >>
rlabel locali s 1826 276 1854 304 4 Clk_Out
port 1 nsew
rlabel metal1 s 0 48 0 48 4 GND
port 2 nsew
rlabel locali s 0 278 0 278 4 Clk_In
port 3 nsew
rlabel metal1 s 0 592 0 592 4 VDD
port 4 nsew
<< end >>
