magic
tech sky130B
magscale 1 2
timestamp 1662180122
<< nwell >>
rect 960 -1180 2385 -750
<< pwell >>
rect 974 -1314 1196 -1224
rect 1594 -1304 1816 -1224
rect 2134 -1304 2366 -1224
rect 1594 -1314 2366 -1304
rect 974 -1476 2366 -1314
rect 1304 -1716 1456 -1476
rect 1844 -1696 2096 -1476
<< nmos >>
rect 1330 -1620 1420 -1420
rect 2230 -1450 2260 -1250
<< pmos >>
rect 2220 -1110 2260 -910
<< pmoslvt >>
rect 1070 -1060 1270 -860
rect 1520 -1060 1720 -860
rect 1930 -1060 2020 -860
<< nmoslvt >>
rect 1070 -1450 1100 -1250
rect 1690 -1450 1720 -1250
rect 1870 -1600 2070 -1400
<< ndiff >>
rect 1000 -1299 1070 -1250
rect 1000 -1333 1013 -1299
rect 1047 -1333 1070 -1299
rect 1000 -1367 1070 -1333
rect 1000 -1401 1013 -1367
rect 1047 -1401 1070 -1367
rect 1000 -1450 1070 -1401
rect 1100 -1299 1170 -1250
rect 1100 -1333 1123 -1299
rect 1157 -1333 1170 -1299
rect 1100 -1367 1170 -1333
rect 1620 -1299 1690 -1250
rect 1620 -1333 1633 -1299
rect 1667 -1333 1690 -1299
rect 1100 -1401 1123 -1367
rect 1157 -1401 1170 -1367
rect 1100 -1450 1170 -1401
rect 1330 -1358 1420 -1340
rect 1330 -1392 1358 -1358
rect 1392 -1392 1420 -1358
rect 1330 -1420 1420 -1392
rect 1620 -1367 1690 -1333
rect 1620 -1401 1633 -1367
rect 1667 -1401 1690 -1367
rect 1620 -1450 1690 -1401
rect 1720 -1299 1790 -1250
rect 1720 -1333 1743 -1299
rect 1777 -1333 1790 -1299
rect 2160 -1299 2230 -1250
rect 1720 -1367 1790 -1333
rect 1720 -1401 1743 -1367
rect 1777 -1401 1790 -1367
rect 1870 -1343 2070 -1330
rect 1870 -1377 1919 -1343
rect 1953 -1377 1987 -1343
rect 2021 -1377 2070 -1343
rect 1870 -1400 2070 -1377
rect 2160 -1333 2173 -1299
rect 2207 -1333 2230 -1299
rect 2160 -1367 2230 -1333
rect 1720 -1450 1790 -1401
rect 2160 -1401 2173 -1367
rect 2207 -1401 2230 -1367
rect 2160 -1450 2230 -1401
rect 2260 -1299 2340 -1250
rect 2260 -1333 2288 -1299
rect 2322 -1333 2340 -1299
rect 2260 -1367 2340 -1333
rect 2260 -1401 2288 -1367
rect 2322 -1401 2340 -1367
rect 2260 -1450 2340 -1401
rect 1330 -1640 1420 -1620
rect 1870 -1623 2070 -1600
rect 1330 -1643 1430 -1640
rect 1330 -1677 1373 -1643
rect 1407 -1677 1430 -1643
rect 1870 -1657 1924 -1623
rect 1958 -1657 1992 -1623
rect 2026 -1657 2070 -1623
rect 1870 -1670 2070 -1657
rect 1330 -1690 1430 -1677
<< pdiff >>
rect 1000 -909 1070 -860
rect 1000 -943 1013 -909
rect 1047 -943 1070 -909
rect 1000 -977 1070 -943
rect 1000 -1011 1013 -977
rect 1047 -1011 1070 -977
rect 1000 -1060 1070 -1011
rect 1270 -909 1350 -860
rect 1450 -909 1520 -860
rect 1270 -943 1293 -909
rect 1327 -943 1350 -909
rect 1450 -943 1471 -909
rect 1505 -943 1520 -909
rect 1270 -977 1350 -943
rect 1450 -977 1520 -943
rect 1270 -1011 1293 -977
rect 1327 -1011 1350 -977
rect 1450 -1011 1471 -977
rect 1505 -1011 1520 -977
rect 1270 -1060 1350 -1011
rect 1450 -1060 1520 -1011
rect 1720 -909 1790 -860
rect 1720 -943 1743 -909
rect 1777 -943 1790 -909
rect 1720 -977 1790 -943
rect 1720 -1011 1743 -977
rect 1777 -1011 1790 -977
rect 1720 -1060 1790 -1011
rect 1860 -909 1930 -860
rect 1860 -943 1873 -909
rect 1907 -943 1930 -909
rect 1860 -977 1930 -943
rect 1860 -1011 1873 -977
rect 1907 -1011 1930 -977
rect 1860 -1060 1930 -1011
rect 2020 -909 2090 -860
rect 2020 -943 2043 -909
rect 2077 -943 2090 -909
rect 2020 -977 2090 -943
rect 2020 -1011 2043 -977
rect 2077 -1011 2090 -977
rect 2020 -1060 2090 -1011
rect 2150 -959 2220 -910
rect 2150 -993 2166 -959
rect 2200 -993 2220 -959
rect 2150 -1027 2220 -993
rect 2150 -1061 2166 -1027
rect 2200 -1061 2220 -1027
rect 2150 -1110 2220 -1061
rect 2260 -959 2330 -910
rect 2260 -993 2283 -959
rect 2317 -993 2330 -959
rect 2260 -1027 2330 -993
rect 2260 -1061 2283 -1027
rect 2317 -1061 2330 -1027
rect 2260 -1110 2330 -1061
<< ndiffc >>
rect 1013 -1333 1047 -1299
rect 1013 -1401 1047 -1367
rect 1123 -1333 1157 -1299
rect 1633 -1333 1667 -1299
rect 1123 -1401 1157 -1367
rect 1358 -1392 1392 -1358
rect 1633 -1401 1667 -1367
rect 1743 -1333 1777 -1299
rect 1743 -1401 1777 -1367
rect 1919 -1377 1953 -1343
rect 1987 -1377 2021 -1343
rect 2173 -1333 2207 -1299
rect 2173 -1401 2207 -1367
rect 2288 -1333 2322 -1299
rect 2288 -1401 2322 -1367
rect 1373 -1677 1407 -1643
rect 1924 -1657 1958 -1623
rect 1992 -1657 2026 -1623
<< pdiffc >>
rect 1013 -943 1047 -909
rect 1013 -1011 1047 -977
rect 1293 -943 1327 -909
rect 1471 -943 1505 -909
rect 1293 -1011 1327 -977
rect 1471 -1011 1505 -977
rect 1743 -943 1777 -909
rect 1743 -1011 1777 -977
rect 1873 -943 1907 -909
rect 1873 -1011 1907 -977
rect 2043 -943 2077 -909
rect 2043 -1011 2077 -977
rect 2166 -993 2200 -959
rect 2166 -1061 2200 -1027
rect 2283 -993 2317 -959
rect 2283 -1061 2317 -1027
<< psubdiff >>
rect 490 -1920 650 -1890
rect 490 -2130 530 -1920
rect 630 -2130 650 -1920
rect 490 -2160 650 -2130
<< nsubdiff >>
rect 1350 -909 1450 -860
rect 1350 -943 1383 -909
rect 1417 -943 1450 -909
rect 1350 -977 1450 -943
rect 1350 -1011 1383 -977
rect 1417 -1011 1450 -977
rect 1350 -1060 1450 -1011
<< psubdiffcont >>
rect 530 -2130 630 -1920
<< nsubdiffcont >>
rect 1383 -943 1417 -909
rect 1383 -1011 1417 -977
<< poly >>
rect 1070 -860 1270 -830
rect 1520 -860 1720 -830
rect 1930 -860 2020 -830
rect 2220 -910 2260 -880
rect 1070 -1090 1270 -1060
rect 1520 -1090 1720 -1060
rect 1930 -1090 2020 -1060
rect 1070 -1123 1150 -1090
rect 1070 -1157 1093 -1123
rect 1127 -1157 1150 -1123
rect 1235 -1130 1550 -1090
rect 1930 -1107 1980 -1090
rect 1918 -1123 1980 -1107
rect 1680 -1143 1720 -1140
rect 1070 -1170 1150 -1157
rect 1617 -1153 1720 -1143
rect 1617 -1187 1633 -1153
rect 1667 -1187 1720 -1153
rect 1918 -1157 1928 -1123
rect 1962 -1157 1980 -1123
rect 2220 -1150 2260 -1110
rect 1918 -1170 1980 -1157
rect 1918 -1173 1972 -1170
rect 1617 -1197 1720 -1187
rect 1680 -1200 1720 -1197
rect 1070 -1250 1100 -1220
rect 1690 -1250 1720 -1200
rect 2027 -1193 2093 -1183
rect 2027 -1227 2043 -1193
rect 2077 -1195 2093 -1193
rect 2230 -1195 2260 -1150
rect 2077 -1225 2260 -1195
rect 2077 -1227 2093 -1225
rect 2027 -1237 2093 -1227
rect 2230 -1250 2260 -1225
rect 1250 -1440 1330 -1420
rect 1070 -1497 1100 -1450
rect 1240 -1489 1330 -1440
rect 1058 -1513 1112 -1497
rect 1058 -1547 1068 -1513
rect 1102 -1547 1112 -1513
rect 1058 -1563 1112 -1547
rect 1240 -1523 1253 -1489
rect 1287 -1523 1330 -1489
rect 1240 -1557 1330 -1523
rect 1240 -1591 1253 -1557
rect 1287 -1591 1330 -1557
rect 1240 -1620 1330 -1591
rect 1420 -1620 1460 -1420
rect 1690 -1480 1720 -1450
rect 1840 -1520 1870 -1400
rect 1770 -1548 1870 -1520
rect 1770 -1582 1793 -1548
rect 1827 -1582 1870 -1548
rect 1770 -1600 1870 -1582
rect 2070 -1600 2100 -1400
rect 2230 -1500 2260 -1450
rect 1770 -1610 1840 -1600
<< polycont >>
rect 1093 -1157 1127 -1123
rect 1633 -1187 1667 -1153
rect 1928 -1157 1962 -1123
rect 2043 -1227 2077 -1193
rect 1068 -1547 1102 -1513
rect 1253 -1523 1287 -1489
rect 1253 -1591 1287 -1557
rect 1793 -1582 1827 -1548
<< locali >>
rect 1350 -740 1450 -730
rect 1100 -758 2270 -740
rect 1100 -792 1179 -758
rect 1213 -792 1251 -758
rect 1285 -792 1323 -758
rect 1357 -792 1395 -758
rect 1429 -792 1467 -758
rect 1501 -792 1539 -758
rect 1573 -792 1611 -758
rect 1645 -792 1683 -758
rect 1717 -792 1755 -758
rect 1789 -792 1827 -758
rect 1861 -792 1899 -758
rect 1933 -792 1971 -758
rect 2005 -792 2043 -758
rect 2077 -792 2115 -758
rect 2149 -792 2187 -758
rect 2221 -792 2270 -758
rect 1100 -810 2270 -792
rect 1350 -860 1450 -810
rect 1000 -909 1050 -860
rect 1000 -943 1013 -909
rect 1047 -943 1050 -909
rect 1000 -977 1050 -943
rect 1000 -1011 1013 -977
rect 1047 -1011 1050 -977
rect 1000 -1123 1050 -1011
rect 1290 -909 1510 -860
rect 1290 -943 1293 -909
rect 1327 -943 1383 -909
rect 1417 -943 1471 -909
rect 1505 -943 1510 -909
rect 1290 -977 1510 -943
rect 1290 -1011 1293 -977
rect 1327 -1011 1383 -977
rect 1417 -1011 1471 -977
rect 1505 -1011 1510 -977
rect 1290 -1060 1510 -1011
rect 1740 -909 1790 -860
rect 1740 -943 1743 -909
rect 1777 -943 1790 -909
rect 1740 -977 1790 -943
rect 1740 -1011 1743 -977
rect 1777 -1011 1790 -977
rect 800 -1500 870 -1130
rect 1000 -1157 1093 -1123
rect 1127 -1157 1143 -1123
rect 1740 -1130 1790 -1011
rect 1860 -909 1910 -810
rect 1860 -943 1873 -909
rect 1907 -943 1910 -909
rect 1860 -977 1910 -943
rect 1860 -1011 1873 -977
rect 1907 -1011 1910 -977
rect 1860 -1060 1910 -1011
rect 2030 -909 2090 -860
rect 2030 -943 2043 -909
rect 2077 -943 2090 -909
rect 2160 -910 2200 -810
rect 2030 -977 2090 -943
rect 2030 -1011 2043 -977
rect 2077 -1011 2090 -977
rect 2030 -1060 2090 -1011
rect 1912 -1130 1928 -1123
rect 1633 -1153 1667 -1137
rect 1000 -1299 1050 -1157
rect 1740 -1157 1928 -1130
rect 1962 -1130 1978 -1123
rect 1962 -1157 1980 -1130
rect 1740 -1170 1980 -1157
rect 1000 -1333 1013 -1299
rect 1047 -1333 1050 -1299
rect 1000 -1367 1050 -1333
rect 1000 -1401 1013 -1367
rect 1047 -1401 1050 -1367
rect 1000 -1450 1050 -1401
rect 1120 -1299 1170 -1250
rect 1120 -1333 1123 -1299
rect 1157 -1333 1170 -1299
rect 1120 -1340 1170 -1333
rect 1620 -1299 1670 -1250
rect 1620 -1333 1633 -1299
rect 1667 -1333 1670 -1299
rect 1620 -1340 1670 -1333
rect 1120 -1358 1670 -1340
rect 1120 -1367 1358 -1358
rect 1120 -1401 1123 -1367
rect 1157 -1392 1358 -1367
rect 1392 -1367 1670 -1358
rect 1392 -1392 1633 -1367
rect 1157 -1400 1633 -1392
rect 1157 -1401 1170 -1400
rect 1120 -1450 1170 -1401
rect 1620 -1401 1633 -1400
rect 1667 -1401 1670 -1367
rect 1240 -1468 1310 -1440
rect 1620 -1450 1670 -1401
rect 1740 -1299 1790 -1170
rect 2040 -1193 2090 -1060
rect 2150 -959 2200 -910
rect 2150 -993 2166 -959
rect 2150 -1027 2200 -993
rect 2150 -1061 2166 -1027
rect 2150 -1110 2200 -1061
rect 2280 -959 2340 -910
rect 2280 -993 2283 -959
rect 2317 -993 2340 -959
rect 2280 -1027 2340 -993
rect 2280 -1061 2283 -1027
rect 2317 -1061 2340 -1027
rect 2040 -1227 2043 -1193
rect 2077 -1227 2090 -1193
rect 2040 -1290 2090 -1227
rect 2280 -1203 2340 -1061
rect 2280 -1237 2293 -1203
rect 2327 -1237 2340 -1203
rect 1740 -1333 1743 -1299
rect 1777 -1333 1790 -1299
rect 1740 -1367 1790 -1333
rect 1740 -1401 1743 -1367
rect 1777 -1401 1790 -1367
rect 1870 -1320 2090 -1290
rect 2150 -1299 2210 -1250
rect 1870 -1343 2070 -1320
rect 1870 -1377 1919 -1343
rect 1953 -1377 1987 -1343
rect 2021 -1377 2070 -1343
rect 1870 -1380 2070 -1377
rect 2150 -1333 2173 -1299
rect 2207 -1333 2210 -1299
rect 2150 -1367 2210 -1333
rect 1740 -1450 1790 -1401
rect 2150 -1401 2173 -1367
rect 2207 -1401 2210 -1367
rect 800 -1513 1120 -1500
rect 800 -1547 1068 -1513
rect 1102 -1547 1120 -1513
rect 800 -1570 1120 -1547
rect 1240 -1523 1253 -1468
rect 1287 -1523 1310 -1468
rect 1780 -1520 1840 -1510
rect 1240 -1557 1310 -1523
rect 1240 -1591 1253 -1557
rect 1287 -1591 1310 -1557
rect 1240 -1620 1310 -1591
rect 1770 -1538 1840 -1520
rect 1770 -1572 1788 -1538
rect 1822 -1548 1840 -1538
rect 1770 -1582 1793 -1572
rect 1827 -1582 1840 -1548
rect 1770 -1610 1840 -1582
rect 1880 -1623 2070 -1610
rect 1350 -1643 1500 -1640
rect 1350 -1677 1372 -1643
rect 1407 -1677 1444 -1643
rect 1478 -1677 1500 -1643
rect 1350 -1690 1500 -1677
rect 1880 -1657 1924 -1623
rect 1958 -1643 1992 -1623
rect 2026 -1640 2070 -1623
rect 2026 -1643 2080 -1640
rect 1961 -1657 1992 -1643
rect 1880 -1677 1927 -1657
rect 1961 -1677 1999 -1657
rect 2033 -1677 2080 -1643
rect 1880 -1690 2080 -1677
rect 2150 -1643 2210 -1401
rect 2280 -1299 2340 -1237
rect 2280 -1333 2288 -1299
rect 2322 -1333 2340 -1299
rect 2280 -1367 2340 -1333
rect 2280 -1401 2288 -1367
rect 2322 -1401 2340 -1367
rect 2280 -1450 2340 -1401
rect 2150 -1677 2163 -1643
rect 2197 -1677 2210 -1643
rect 2150 -1690 2210 -1677
rect 490 -1910 650 -1890
rect 490 -2140 510 -1910
rect 640 -2140 650 -1910
rect 770 -1981 810 -1980
rect 764 -2030 813 -1981
rect 490 -2160 650 -2140
rect 770 -2150 810 -2030
rect 1640 -2140 1680 -1970
<< viali >>
rect 1179 -792 1213 -758
rect 1251 -792 1285 -758
rect 1323 -792 1357 -758
rect 1395 -792 1429 -758
rect 1467 -792 1501 -758
rect 1539 -792 1573 -758
rect 1611 -792 1645 -758
rect 1683 -792 1717 -758
rect 1755 -792 1789 -758
rect 1827 -792 1861 -758
rect 1899 -792 1933 -758
rect 1971 -792 2005 -758
rect 2043 -792 2077 -758
rect 2115 -792 2149 -758
rect 2187 -792 2221 -758
rect 1633 -1187 1667 -1178
rect 1633 -1212 1667 -1187
rect 2293 -1237 2327 -1203
rect 1068 -1547 1102 -1513
rect 1253 -1489 1287 -1468
rect 1253 -1502 1287 -1489
rect 1788 -1548 1822 -1538
rect 1788 -1572 1793 -1548
rect 1793 -1572 1822 -1548
rect 1372 -1677 1373 -1643
rect 1373 -1677 1406 -1643
rect 1444 -1677 1478 -1643
rect 1927 -1657 1958 -1643
rect 1958 -1657 1961 -1643
rect 1999 -1657 2026 -1643
rect 2026 -1657 2033 -1643
rect 1927 -1677 1961 -1657
rect 1999 -1677 2033 -1657
rect 2163 -1677 2197 -1643
rect 510 -1920 640 -1910
rect 510 -2130 530 -1920
rect 530 -2130 630 -1920
rect 630 -2130 640 -1920
rect 510 -2140 640 -2130
<< metal1 >>
rect 760 -758 2290 -730
rect 760 -792 1179 -758
rect 1213 -792 1251 -758
rect 1285 -792 1323 -758
rect 1357 -792 1395 -758
rect 1429 -792 1467 -758
rect 1501 -792 1539 -758
rect 1573 -792 1611 -758
rect 1645 -792 1683 -758
rect 1717 -792 1755 -758
rect 1789 -792 1827 -758
rect 1861 -792 1899 -758
rect 1933 -792 1971 -758
rect 2005 -792 2043 -758
rect 2077 -792 2115 -758
rect 2149 -792 2187 -758
rect 2221 -770 2290 -758
rect 2221 -792 2500 -770
rect 760 -830 2500 -792
rect 1624 -1169 1676 -1163
rect 2274 -1180 2346 -1178
rect 1624 -1227 1676 -1221
rect 2270 -1199 2390 -1180
rect 2270 -1203 2314 -1199
rect 2270 -1237 2293 -1203
rect 2270 -1251 2314 -1237
rect 2366 -1251 2390 -1199
rect 2270 -1270 2390 -1251
rect 660 -1410 2500 -1350
rect 1230 -1468 1310 -1440
rect 1230 -1488 1253 -1468
rect 1214 -1494 1253 -1488
rect 1062 -1504 1108 -1501
rect 1287 -1502 1310 -1468
rect 1053 -1556 1059 -1504
rect 1111 -1556 1117 -1504
rect 1266 -1530 1310 -1502
rect 1760 -1510 1790 -1410
rect 1760 -1520 1840 -1510
rect 1214 -1552 1266 -1546
rect 1760 -1538 1850 -1520
rect 1062 -1559 1108 -1556
rect 1760 -1572 1788 -1538
rect 1822 -1572 1850 -1538
rect 1760 -1590 1850 -1572
rect 660 -1625 705 -1615
rect 660 -1643 2330 -1625
rect 660 -1677 1372 -1643
rect 1406 -1677 1444 -1643
rect 1478 -1677 1927 -1643
rect 1961 -1677 1999 -1643
rect 2033 -1677 2163 -1643
rect 2197 -1677 2330 -1643
rect 660 -1695 2330 -1677
rect 660 -1830 705 -1695
rect 450 -1910 705 -1830
rect 450 -2140 510 -1910
rect 640 -2140 705 -1910
rect 450 -2180 705 -2140
rect 660 -2360 705 -2180
<< via1 >>
rect 1624 -1178 1676 -1169
rect 1624 -1212 1633 -1178
rect 1633 -1212 1667 -1178
rect 1667 -1212 1676 -1178
rect 1624 -1221 1676 -1212
rect 2314 -1203 2366 -1199
rect 2314 -1237 2327 -1203
rect 2327 -1237 2366 -1203
rect 2314 -1251 2366 -1237
rect 1214 -1502 1253 -1494
rect 1253 -1502 1266 -1494
rect 1059 -1513 1111 -1504
rect 1059 -1547 1068 -1513
rect 1068 -1547 1102 -1513
rect 1102 -1547 1111 -1513
rect 1059 -1556 1111 -1547
rect 1214 -1546 1266 -1502
<< metal2 >>
rect 939 -885 969 -665
rect 939 -915 970 -885
rect 939 -1735 969 -915
rect 1059 -1504 1111 -1498
rect 1059 -1562 1111 -1556
rect 1140 -1630 1180 -720
rect 1210 -1492 1270 -1481
rect 1210 -1494 1212 -1492
rect 1268 -1494 1270 -1492
rect 1208 -1546 1212 -1494
rect 1268 -1546 1272 -1494
rect 1210 -1548 1212 -1546
rect 1268 -1548 1270 -1546
rect 1210 -1559 1270 -1548
rect 1104 -1670 1180 -1630
rect 1104 -1730 1144 -1670
rect 1374 -1735 1404 -720
rect 1539 -1730 1579 -720
rect 1610 -922 1690 -901
rect 1610 -978 1622 -922
rect 1678 -978 1690 -922
rect 1610 -1169 1690 -978
rect 1610 -1221 1624 -1169
rect 1676 -1221 1690 -1169
rect 1610 -1240 1690 -1221
rect 1809 -1725 1839 -720
rect 1974 -1740 2014 -720
rect 2244 -805 2274 -695
rect 2236 -806 2274 -805
rect 2205 -835 2274 -806
rect 2205 -1345 2235 -835
rect 2409 -1040 2449 -720
rect 2410 -1060 2449 -1040
rect 2410 -1100 2500 -1060
rect 2300 -1199 2390 -1180
rect 2300 -1200 2314 -1199
rect 2366 -1200 2390 -1199
rect 2300 -1260 2310 -1200
rect 2370 -1260 2390 -1200
rect 2300 -1270 2390 -1260
rect 2470 -1310 2500 -1100
rect 2205 -1375 2274 -1345
rect 2244 -1735 2274 -1375
rect 2409 -1350 2500 -1310
rect 2409 -1700 2449 -1350
<< via2 >>
rect 1212 -1494 1268 -1492
rect 1212 -1546 1214 -1494
rect 1214 -1546 1266 -1494
rect 1266 -1546 1268 -1494
rect 1212 -1548 1268 -1546
rect 1622 -978 1678 -922
rect 2310 -1251 2314 -1200
rect 2314 -1251 2366 -1200
rect 2366 -1251 2370 -1200
rect 2310 -1260 2370 -1251
<< metal3 >>
rect 920 -922 2620 -900
rect 920 -960 1622 -922
rect 1605 -978 1622 -960
rect 1678 -960 2620 -922
rect 1678 -978 1695 -960
rect 1605 -995 1695 -978
rect 920 -1130 2630 -1070
rect 1210 -1485 1270 -1130
rect 2300 -1200 2390 -1190
rect 2300 -1260 2310 -1200
rect 2370 -1260 2390 -1200
rect 2300 -1445 2390 -1260
rect 1205 -1492 1275 -1485
rect 1205 -1548 1212 -1492
rect 1268 -1548 1275 -1492
rect 2300 -1535 2545 -1445
rect 1205 -1555 1275 -1548
rect 2455 -1795 2545 -1535
rect 540 -2320 2500 -2260
<< metal4 >>
rect 814 -1750 874 -680
rect 1004 -1740 1064 -680
rect 1249 -1740 1309 -720
rect 1439 -1740 1499 -720
rect 1684 -1740 1744 -720
rect 1874 -1740 1934 -720
rect 2119 -1740 2179 -720
rect 2309 -1740 2369 -720
use 8bit_dram  8bit_dram_0
timestamp 1662167647
transform -1 0 2469 0 -1 -1700
box -70 -20 1745 780
<< labels >>
rlabel locali 830 -1150 830 -1150 1 V_IN
port 1 n
rlabel metal1 680 -1380 680 -1380 1 BIAS2
port 2 n
rlabel metal1 730 -1660 730 -1660 1 GND
port 3 n
rlabel metal3 2530 -1100 2530 -1100 1 BIAS1
port 4 n
rlabel metal1 810 -770 810 -770 1 VDD
port 5 n
rlabel metal3 2530 -930 2530 -930 1 V_RAMP
port 6 n
rlabel metal4 2340 -730 2340 -730 1 GRAY_INx1x
port 7 n
rlabel metal2 2430 -730 2430 -730 1 GRAY_INx0x
port 8 n
rlabel metal2 2260 -710 2260 -710 1 OUTx1x
port 9 n
rlabel metal4 2150 -720 2150 -720 1 OUTx0x
port 10 n
rlabel metal2 1990 -720 1990 -720 1 GRAY_INx2x
port 11 n
rlabel metal4 1900 -720 1900 -720 1 GRAY_INx3x
port 12 n
rlabel metal2 1820 -720 1820 -720 1 OUTx3x
port 13 n
rlabel metal4 1710 -720 1710 -720 1 OUTx2x
port 14 n
rlabel metal2 1560 -720 1560 -720 1 GRAY_INx4x
port 15 n
rlabel metal4 1470 -720 1470 -720 1 GRAY_INx5x
port 16 n
rlabel metal2 1390 -720 1390 -720 1 OUTx5x
port 17 n
rlabel metal4 1280 -720 1280 -720 1 OUTx4x
port 18 n
rlabel metal2 1160 -720 1160 -720 1 GRAY_INx6x
port 19 n
rlabel metal4 1030 -700 1030 -700 1 GRAY_INx7x
port 20 n
rlabel metal2 950 -690 950 -690 1 OUTx7x
port 21 n
rlabel metal4 840 -700 840 -700 1 OUTx6x
port 22 n
rlabel metal3 570 -2290 570 -2290 1 READ
port 23 n
<< end >>
