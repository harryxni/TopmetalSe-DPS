** sch_path: /home/hni/topmetal_dps/xschem/testbench/sens_amp_tb.sch
**.subckt sens_amp_tb
x5 OUT VREF TEST SA_IREF sens_amp
I8 VDD SA_IREF 200n
XM7 GND SA_IREF SA_IREF GND sky130_fd_pr__nfet_01v8_lvt L=1 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
V10 VREF GND 400m
V8 VDD GND 1.8
V1 TEST GND PULSE(0 800m 10u 0.01u 0.01u 10u)
**** begin user architecture code

** opencircuitdesign pdks install
.lib /opt/OpenICEDA/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends

* expanding   symbol:  sens_amp.sym # of pins=4
** sym_path: /home/hni/topmetal_dps/xschem/sens_amp.sym
** sch_path: /home/hni/topmetal_dps/xschem/sens_amp.sch
.subckt sens_amp  OUT REF V_IN SA_IREF
*.ipin REF
*.ipin V_IN
*.opin OUT
*.ipin SA_IREF
X0 GN GN VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=3.5e+11p pd=2.7e+06u as=1.8e+12p ps=1.22e+07u w=1e+06u l=500000u
X1 net1 V_IN net2 GND sky130_fd_pr__nfet_01v8_lvt ad=1.4e+12p pd=8.7e+06u as=1.775e+12p ps=1.05e+07u w=4e+06u l=150000u
X2 net2 REF GN GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+12p ps=9.1e+06u w=4e+06u l=150000u
X3 net1 GN VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=3.5e+11p pd=2.7e+06u as=0p ps=0u w=1e+06u l=500000u
X4 net2 SA_IREF GND GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=6e+11p ps=4.7e+06u w=500000u l=1e+06u
X5 OUT net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.05e+12p pd=6.7e+06u as=0p ps=0u w=3e+06u l=350000u
X6 OUT net1 GND GND sky130_fd_pr__nfet_01v8_lvt ad=3.5e+11p pd=2.7e+06u as=0p ps=0u w=1e+06u l=150000u




.ends

.GLOBAL GND
.GLOBAL VDD
**** begin user architecture code


.options gmin=10e-20
.control
save all

*dc v2 0 1.8 0.05
*plot v(test)
tran 1u 200u

write sim_dpspixel_tb.raw
.endc


**** end user architecture code
.end
