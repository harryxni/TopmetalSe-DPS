magic
tech sky130B
magscale 1 2
timestamp 1607746020
<< locali >>
rect 14197 2839 14231 3145
rect 36829 2907 36863 3145
rect 42165 2839 42199 3009
rect 45845 2907 45879 3077
rect 12633 1411 12667 1513
<< viali >>
rect 14197 3145 14231 3179
rect 2789 3009 2823 3043
rect 3617 3009 3651 3043
rect 3893 3009 3927 3043
rect 4537 3009 4571 3043
rect 4905 3009 4939 3043
rect 5825 3009 5859 3043
rect 6377 3009 6411 3043
rect 7205 3009 7239 3043
rect 8493 3009 8527 3043
rect 8769 3009 8803 3043
rect 9689 3009 9723 3043
rect 10057 3009 10091 3043
rect 11713 3009 11747 3043
rect 12909 3009 12943 3043
rect 13277 3009 13311 3043
rect 3065 2941 3099 2975
rect 3341 2941 3375 2975
rect 5181 2941 5215 2975
rect 6653 2941 6687 2975
rect 7481 2941 7515 2975
rect 9045 2941 9079 2975
rect 10333 2941 10367 2975
rect 11345 2941 11379 2975
rect 13645 2941 13679 2975
rect 1961 2873 1995 2907
rect 7941 2873 7975 2907
rect 9321 2873 9355 2907
rect 10609 2873 10643 2907
rect 12265 2873 12299 2907
rect 36829 3145 36863 3179
rect 15393 3009 15427 3043
rect 15761 3009 15795 3043
rect 17417 3009 17451 3043
rect 17693 3009 17727 3043
rect 19533 3009 19567 3043
rect 20177 3009 20211 3043
rect 21097 3009 21131 3043
rect 21465 3009 21499 3043
rect 22109 3009 22143 3043
rect 22661 3009 22695 3043
rect 22937 3009 22971 3043
rect 24317 3009 24351 3043
rect 25605 3009 25639 3043
rect 28181 3009 28215 3043
rect 28457 3009 28491 3043
rect 31585 3009 31619 3043
rect 31861 3009 31895 3043
rect 32413 3009 32447 3043
rect 32873 3009 32907 3043
rect 33149 3009 33183 3043
rect 33701 3009 33735 3043
rect 34529 3009 34563 3043
rect 35725 3009 35759 3043
rect 36001 3009 36035 3043
rect 14841 2941 14875 2975
rect 16221 2941 16255 2975
rect 16773 2941 16807 2975
rect 19901 2941 19935 2975
rect 21833 2941 21867 2975
rect 23581 2941 23615 2975
rect 32137 2941 32171 2975
rect 33425 2941 33459 2975
rect 35265 2941 35299 2975
rect 45845 3077 45879 3111
rect 37933 3009 37967 3043
rect 40417 3009 40451 3043
rect 40785 3009 40819 3043
rect 41061 3009 41095 3043
rect 42165 3009 42199 3043
rect 42901 3009 42935 3043
rect 43177 3009 43211 3043
rect 43637 3009 43671 3043
rect 44833 3009 44867 3043
rect 45293 3009 45327 3043
rect 38577 2941 38611 2975
rect 41889 2941 41923 2975
rect 14289 2873 14323 2907
rect 15117 2873 15151 2907
rect 17049 2873 17083 2907
rect 18613 2873 18647 2907
rect 18889 2873 18923 2907
rect 20545 2873 20579 2907
rect 22385 2873 22419 2907
rect 23213 2873 23247 2907
rect 28733 2873 28767 2907
rect 30665 2873 30699 2907
rect 34253 2873 34287 2907
rect 34989 2873 35023 2907
rect 36553 2873 36587 2907
rect 36829 2873 36863 2907
rect 36921 2873 36955 2907
rect 38209 2873 38243 2907
rect 40049 2873 40083 2907
rect 44557 2941 44591 2975
rect 47317 3009 47351 3043
rect 47593 3009 47627 3043
rect 48329 3009 48363 3043
rect 49341 3009 49375 3043
rect 49617 3009 49651 3043
rect 50721 3009 50755 3043
rect 50997 3009 51031 3043
rect 52009 3009 52043 3043
rect 53113 3009 53147 3043
rect 53941 3009 53975 3043
rect 54217 3009 54251 3043
rect 55137 3009 55171 3043
rect 56241 3009 56275 3043
rect 56793 3009 56827 3043
rect 57621 3009 57655 3043
rect 46305 2941 46339 2975
rect 48697 2941 48731 2975
rect 49985 2941 50019 2975
rect 51733 2941 51767 2975
rect 52837 2941 52871 2975
rect 54769 2941 54803 2975
rect 55965 2941 55999 2975
rect 57345 2941 57379 2975
rect 42257 2873 42291 2907
rect 43913 2873 43947 2907
rect 45569 2873 45603 2907
rect 45845 2873 45879 2907
rect 46581 2873 46615 2907
rect 48973 2873 49007 2907
rect 50261 2873 50295 2907
rect 51365 2873 51399 2907
rect 52377 2873 52411 2907
rect 53573 2873 53607 2907
rect 54493 2873 54527 2907
rect 55689 2873 55723 2907
rect 57069 2873 57103 2907
rect 2237 2805 2271 2839
rect 2513 2805 2547 2839
rect 5549 2805 5583 2839
rect 6101 2805 6135 2839
rect 8217 2805 8251 2839
rect 10977 2805 11011 2839
rect 11989 2805 12023 2839
rect 12541 2805 12575 2839
rect 13921 2805 13955 2839
rect 14197 2805 14231 2839
rect 14565 2805 14599 2839
rect 16497 2805 16531 2839
rect 18061 2805 18095 2839
rect 19165 2805 19199 2839
rect 20821 2805 20855 2839
rect 23857 2805 23891 2839
rect 36277 2805 36311 2839
rect 37197 2805 37231 2839
rect 37657 2805 37691 2839
rect 38853 2805 38887 2839
rect 39129 2805 39163 2839
rect 39405 2805 39439 2839
rect 39681 2805 39715 2839
rect 41613 2805 41647 2839
rect 42165 2805 42199 2839
rect 42625 2805 42659 2839
rect 44281 2805 44315 2839
rect 46029 2805 46063 2839
rect 48053 2805 48087 2839
rect 56517 2805 56551 2839
rect 2881 2601 2915 2635
rect 3157 2601 3191 2635
rect 4629 2601 4663 2635
rect 9137 2601 9171 2635
rect 11161 2601 11195 2635
rect 13093 2601 13127 2635
rect 16865 2601 16899 2635
rect 18981 2601 19015 2635
rect 21189 2601 21223 2635
rect 22017 2601 22051 2635
rect 23213 2601 23247 2635
rect 23857 2601 23891 2635
rect 24685 2601 24719 2635
rect 24961 2601 24995 2635
rect 25421 2601 25455 2635
rect 25881 2601 25915 2635
rect 26249 2601 26283 2635
rect 26801 2601 26835 2635
rect 27077 2601 27111 2635
rect 27721 2601 27755 2635
rect 28641 2601 28675 2635
rect 29653 2601 29687 2635
rect 29929 2601 29963 2635
rect 30481 2601 30515 2635
rect 30757 2601 30791 2635
rect 31861 2601 31895 2635
rect 33057 2601 33091 2635
rect 34069 2601 34103 2635
rect 34989 2601 35023 2635
rect 35909 2601 35943 2635
rect 38485 2601 38519 2635
rect 41981 2601 42015 2635
rect 45201 2601 45235 2635
rect 47133 2601 47167 2635
rect 50353 2601 50387 2635
rect 51181 2601 51215 2635
rect 53297 2601 53331 2635
rect 55413 2601 55447 2635
rect 56241 2601 56275 2635
rect 56793 2601 56827 2635
rect 3433 2533 3467 2567
rect 4353 2533 4387 2567
rect 19349 2533 19383 2567
rect 20545 2533 20579 2567
rect 21557 2533 21591 2567
rect 22753 2533 22787 2567
rect 23581 2533 23615 2567
rect 27353 2533 27387 2567
rect 27997 2533 28031 2567
rect 28365 2533 28399 2567
rect 29377 2533 29411 2567
rect 30205 2533 30239 2567
rect 32413 2533 32447 2567
rect 32689 2533 32723 2567
rect 34345 2533 34379 2567
rect 40969 2533 41003 2567
rect 44557 2533 44591 2567
rect 47869 2533 47903 2567
rect 54861 2533 54895 2567
rect 56517 2533 56551 2567
rect 4905 2465 4939 2499
rect 22477 2465 22511 2499
rect 24317 2465 24351 2499
rect 33609 2465 33643 2499
rect 34713 2465 34747 2499
rect 55137 2465 55171 2499
rect 57069 2465 57103 2499
rect 3709 2397 3743 2431
rect 3985 2397 4019 2431
rect 20821 2397 20855 2431
rect 28917 2397 28951 2431
rect 33333 2397 33367 2431
rect 55689 2397 55723 2431
rect 55965 2397 55999 2431
rect 3709 1921 3743 1955
rect 3985 1921 4019 1955
rect 5365 1921 5399 1955
rect 20821 1921 20855 1955
rect 21097 1921 21131 1955
rect 21373 1921 21407 1955
rect 22201 1921 22235 1955
rect 23121 1921 23155 1955
rect 23397 1921 23431 1955
rect 24041 1921 24075 1955
rect 25053 1921 25087 1955
rect 25329 1921 25363 1955
rect 25605 1921 25639 1955
rect 30389 1921 30423 1955
rect 31125 1921 31159 1955
rect 33885 1921 33919 1955
rect 39497 1921 39531 1955
rect 54493 1921 54527 1955
rect 55689 1921 55723 1955
rect 55965 1921 55999 1955
rect 56241 1921 56275 1955
rect 3433 1853 3467 1887
rect 4537 1853 4571 1887
rect 5089 1853 5123 1887
rect 11345 1853 11379 1887
rect 13001 1853 13035 1887
rect 13553 1853 13587 1887
rect 21649 1853 21683 1887
rect 24317 1853 24351 1887
rect 26157 1853 26191 1887
rect 26433 1853 26467 1887
rect 42349 1853 42383 1887
rect 54769 1853 54803 1887
rect 57069 1853 57103 1887
rect 3157 1785 3191 1819
rect 4813 1785 4847 1819
rect 5641 1785 5675 1819
rect 12081 1785 12115 1819
rect 21925 1785 21959 1819
rect 22477 1785 22511 1819
rect 24777 1785 24811 1819
rect 45201 1785 45235 1819
rect 56793 1785 56827 1819
rect 2881 1717 2915 1751
rect 4261 1717 4295 1751
rect 8033 1717 8067 1751
rect 10609 1717 10643 1751
rect 12725 1717 12759 1751
rect 13277 1717 13311 1751
rect 13829 1717 13863 1751
rect 14473 1717 14507 1751
rect 17049 1717 17083 1751
rect 18613 1717 18647 1751
rect 22753 1717 22787 1751
rect 25881 1717 25915 1751
rect 27997 1717 28031 1751
rect 37933 1717 37967 1751
rect 41153 1717 41187 1751
rect 43177 1717 43211 1751
rect 48329 1717 48363 1751
rect 49985 1717 50019 1751
rect 55229 1717 55263 1751
rect 56517 1717 56551 1751
rect 57621 1717 57655 1751
rect 2881 1513 2915 1547
rect 4629 1513 4663 1547
rect 7849 1513 7883 1547
rect 9321 1513 9355 1547
rect 11253 1513 11287 1547
rect 12357 1513 12391 1547
rect 12633 1513 12667 1547
rect 13461 1513 13495 1547
rect 14289 1513 14323 1547
rect 19717 1513 19751 1547
rect 20913 1513 20947 1547
rect 22937 1513 22971 1547
rect 24317 1513 24351 1547
rect 24869 1513 24903 1547
rect 25145 1513 25179 1547
rect 27721 1513 27755 1547
rect 28365 1513 28399 1547
rect 29193 1513 29227 1547
rect 30665 1513 30699 1547
rect 31585 1513 31619 1547
rect 32229 1513 32263 1547
rect 34161 1513 34195 1547
rect 34437 1513 34471 1547
rect 34805 1513 34839 1547
rect 35081 1513 35115 1547
rect 35725 1513 35759 1547
rect 36829 1513 36863 1547
rect 37381 1513 37415 1547
rect 39221 1513 39255 1547
rect 41797 1513 41831 1547
rect 43729 1513 43763 1547
rect 44925 1513 44959 1547
rect 46765 1513 46799 1547
rect 48145 1513 48179 1547
rect 49341 1513 49375 1547
rect 50169 1513 50203 1547
rect 51365 1513 51399 1547
rect 52193 1513 52227 1547
rect 55689 1513 55723 1547
rect 55965 1513 55999 1547
rect 56793 1513 56827 1547
rect 2053 1445 2087 1479
rect 3433 1445 3467 1479
rect 3985 1445 4019 1479
rect 5641 1445 5675 1479
rect 6285 1445 6319 1479
rect 7205 1445 7239 1479
rect 8217 1445 8251 1479
rect 9045 1445 9079 1479
rect 10241 1445 10275 1479
rect 11897 1445 11931 1479
rect 13185 1445 13219 1479
rect 16957 1445 16991 1479
rect 18061 1445 18095 1479
rect 19073 1445 19107 1479
rect 20637 1445 20671 1479
rect 21465 1445 21499 1479
rect 23397 1445 23431 1479
rect 26065 1445 26099 1479
rect 26341 1445 26375 1479
rect 26617 1445 26651 1479
rect 27169 1445 27203 1479
rect 28641 1445 28675 1479
rect 30941 1445 30975 1479
rect 31217 1445 31251 1479
rect 32505 1445 32539 1479
rect 33885 1445 33919 1479
rect 35357 1445 35391 1479
rect 37657 1445 37691 1479
rect 37933 1445 37967 1479
rect 40233 1445 40267 1479
rect 40877 1445 40911 1479
rect 42165 1445 42199 1479
rect 42993 1445 43027 1479
rect 45201 1445 45235 1479
rect 47133 1445 47167 1479
rect 48421 1445 48455 1479
rect 50445 1445 50479 1479
rect 51089 1445 51123 1479
rect 52469 1445 52503 1479
rect 53113 1445 53147 1479
rect 53757 1445 53791 1479
rect 54401 1445 54435 1479
rect 55321 1445 55355 1479
rect 57345 1445 57379 1479
rect 57897 1445 57931 1479
rect 2329 1377 2363 1411
rect 2605 1377 2639 1411
rect 3157 1377 3191 1411
rect 4353 1377 4387 1411
rect 4905 1377 4939 1411
rect 5365 1377 5399 1411
rect 6009 1377 6043 1411
rect 6653 1377 6687 1411
rect 7573 1377 7607 1411
rect 8769 1377 8803 1411
rect 9597 1377 9631 1411
rect 10977 1377 11011 1411
rect 11529 1377 11563 1411
rect 12633 1377 12667 1411
rect 12909 1377 12943 1411
rect 13737 1377 13771 1411
rect 14013 1377 14047 1411
rect 14657 1377 14691 1411
rect 15025 1377 15059 1411
rect 15301 1377 15335 1411
rect 15761 1377 15795 1411
rect 16037 1377 16071 1411
rect 16405 1377 16439 1411
rect 16681 1377 16715 1411
rect 17325 1377 17359 1411
rect 17785 1377 17819 1411
rect 19441 1377 19475 1411
rect 20085 1377 20119 1411
rect 20361 1377 20395 1411
rect 21925 1377 21959 1411
rect 22569 1377 22603 1411
rect 24593 1377 24627 1411
rect 25421 1377 25455 1411
rect 25789 1377 25823 1411
rect 27997 1377 28031 1411
rect 30297 1377 30331 1411
rect 32873 1377 32907 1411
rect 33241 1377 33275 1411
rect 33609 1377 33643 1411
rect 36001 1377 36035 1411
rect 37105 1377 37139 1411
rect 38577 1377 38611 1411
rect 39865 1377 39899 1411
rect 40509 1377 40543 1411
rect 41521 1377 41555 1411
rect 42533 1377 42567 1411
rect 44373 1377 44407 1411
rect 44649 1377 44683 1411
rect 45753 1377 45787 1411
rect 46489 1377 46523 1411
rect 47777 1377 47811 1411
rect 48697 1377 48731 1411
rect 49617 1377 49651 1411
rect 50813 1377 50847 1411
rect 51641 1377 51675 1411
rect 53389 1377 53423 1411
rect 54033 1377 54067 1411
rect 54677 1377 54711 1411
rect 54953 1377 54987 1411
rect 56241 1377 56275 1411
rect 56517 1377 56551 1411
rect 3709 1309 3743 1343
rect 8493 1309 8527 1343
rect 10517 1309 10551 1343
rect 18613 1309 18647 1343
rect 22293 1309 22327 1343
rect 23765 1309 23799 1343
rect 27445 1309 27479 1343
rect 28917 1309 28951 1343
rect 29561 1309 29595 1343
rect 30021 1309 30055 1343
rect 31861 1309 31895 1343
rect 36461 1309 36495 1343
rect 38209 1309 38243 1343
rect 38945 1309 38979 1343
rect 39589 1309 39623 1343
rect 43453 1309 43487 1343
rect 45477 1309 45511 1343
rect 46213 1309 46247 1343
rect 47501 1309 47535 1343
rect 48973 1309 49007 1343
rect 52837 1309 52871 1343
rect 57069 1309 57103 1343
rect 57621 1309 57655 1343
<< metal1 >>
rect 16758 3612 16764 3664
rect 16816 3652 16822 3664
rect 18874 3652 18880 3664
rect 16816 3624 18880 3652
rect 16816 3612 16822 3624
rect 18874 3612 18880 3624
rect 18932 3612 18938 3664
rect 31570 3544 31576 3596
rect 31628 3584 31634 3596
rect 35158 3584 35164 3596
rect 31628 3556 35164 3584
rect 31628 3544 31634 3556
rect 35158 3544 35164 3556
rect 35216 3544 35222 3596
rect 15102 3476 15108 3528
rect 15160 3516 15166 3528
rect 16758 3516 16764 3528
rect 15160 3488 16764 3516
rect 15160 3476 15166 3488
rect 16758 3476 16764 3488
rect 16816 3476 16822 3528
rect 33226 3476 33232 3528
rect 33284 3516 33290 3528
rect 35894 3516 35900 3528
rect 33284 3488 35900 3516
rect 33284 3476 33290 3488
rect 35894 3476 35900 3488
rect 35952 3476 35958 3528
rect 19334 3408 19340 3460
rect 19392 3448 19398 3460
rect 22554 3448 22560 3460
rect 19392 3420 22560 3448
rect 19392 3408 19398 3420
rect 22554 3408 22560 3420
rect 22612 3408 22618 3460
rect 33778 3408 33784 3460
rect 33836 3448 33842 3460
rect 36078 3448 36084 3460
rect 33836 3420 36084 3448
rect 33836 3408 33842 3420
rect 36078 3408 36084 3420
rect 36136 3408 36142 3460
rect 36170 3408 36176 3460
rect 36228 3448 36234 3460
rect 36998 3448 37004 3460
rect 36228 3420 37004 3448
rect 36228 3408 36234 3420
rect 36998 3408 37004 3420
rect 37056 3408 37062 3460
rect 37274 3408 37280 3460
rect 37332 3448 37338 3460
rect 38286 3448 38292 3460
rect 37332 3420 38292 3448
rect 37332 3408 37338 3420
rect 38286 3408 38292 3420
rect 38344 3408 38350 3460
rect 38838 3408 38844 3460
rect 38896 3448 38902 3460
rect 40678 3448 40684 3460
rect 38896 3420 40684 3448
rect 38896 3408 38902 3420
rect 40678 3408 40684 3420
rect 40736 3408 40742 3460
rect 19886 3340 19892 3392
rect 19944 3380 19950 3392
rect 22186 3380 22192 3392
rect 19944 3352 22192 3380
rect 19944 3340 19950 3352
rect 22186 3340 22192 3352
rect 22244 3340 22250 3392
rect 34514 3340 34520 3392
rect 34572 3380 34578 3392
rect 35526 3380 35532 3392
rect 34572 3352 35532 3380
rect 34572 3340 34578 3352
rect 35526 3340 35532 3352
rect 35584 3340 35590 3392
rect 36906 3340 36912 3392
rect 36964 3380 36970 3392
rect 38746 3380 38752 3392
rect 36964 3352 38752 3380
rect 36964 3340 36970 3352
rect 38746 3340 38752 3352
rect 38804 3340 38810 3392
rect 39114 3340 39120 3392
rect 39172 3380 39178 3392
rect 40862 3380 40868 3392
rect 39172 3352 40868 3380
rect 39172 3340 39178 3352
rect 40862 3340 40868 3352
rect 40920 3340 40926 3392
rect 42794 3340 42800 3392
rect 42852 3380 42858 3392
rect 43254 3380 43260 3392
rect 42852 3352 43260 3380
rect 42852 3340 42858 3352
rect 43254 3340 43260 3352
rect 43312 3340 43318 3392
rect 44266 3340 44272 3392
rect 44324 3380 44330 3392
rect 45094 3380 45100 3392
rect 44324 3352 45100 3380
rect 44324 3340 44330 3352
rect 45094 3340 45100 3352
rect 45152 3340 45158 3392
rect 1380 3290 58604 3312
rect 1380 3238 3354 3290
rect 3406 3238 19354 3290
rect 19406 3238 35354 3290
rect 35406 3238 51354 3290
rect 51406 3238 58604 3290
rect 1380 3216 58604 3238
rect 842 3136 848 3188
rect 900 3176 906 3188
rect 5074 3176 5080 3188
rect 900 3148 5080 3176
rect 900 3136 906 3148
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 13262 3136 13268 3188
rect 13320 3176 13326 3188
rect 14185 3179 14243 3185
rect 14185 3176 14197 3179
rect 13320 3148 14197 3176
rect 13320 3136 13326 3148
rect 14185 3145 14197 3148
rect 14231 3145 14243 3179
rect 14185 3139 14243 3145
rect 14366 3136 14372 3188
rect 14424 3176 14430 3188
rect 14424 3148 15792 3176
rect 14424 3136 14430 3148
rect 1670 3068 1676 3120
rect 1728 3108 1734 3120
rect 3234 3108 3240 3120
rect 1728 3080 3240 3108
rect 1728 3068 1734 3080
rect 3234 3068 3240 3080
rect 3292 3068 3298 3120
rect 7926 3068 7932 3120
rect 7984 3108 7990 3120
rect 7984 3080 8800 3108
rect 7984 3068 7990 3080
rect 2222 3000 2228 3052
rect 2280 3040 2286 3052
rect 2777 3043 2835 3049
rect 2777 3040 2789 3043
rect 2280 3012 2789 3040
rect 2280 3000 2286 3012
rect 2777 3009 2789 3012
rect 2823 3009 2835 3043
rect 2777 3003 2835 3009
rect 2958 3000 2964 3052
rect 3016 3040 3022 3052
rect 3605 3043 3663 3049
rect 3605 3040 3617 3043
rect 3016 3012 3617 3040
rect 3016 3000 3022 3012
rect 3605 3009 3617 3012
rect 3651 3009 3663 3043
rect 3605 3003 3663 3009
rect 3694 3000 3700 3052
rect 3752 3040 3758 3052
rect 3881 3043 3939 3049
rect 3881 3040 3893 3043
rect 3752 3012 3893 3040
rect 3752 3000 3758 3012
rect 3881 3009 3893 3012
rect 3927 3009 3939 3043
rect 3881 3003 3939 3009
rect 4246 3000 4252 3052
rect 4304 3040 4310 3052
rect 4525 3043 4583 3049
rect 4525 3040 4537 3043
rect 4304 3012 4537 3040
rect 4304 3000 4310 3012
rect 4525 3009 4537 3012
rect 4571 3009 4583 3043
rect 4525 3003 4583 3009
rect 4614 3000 4620 3052
rect 4672 3040 4678 3052
rect 4893 3043 4951 3049
rect 4893 3040 4905 3043
rect 4672 3012 4905 3040
rect 4672 3000 4678 3012
rect 4893 3009 4905 3012
rect 4939 3009 4951 3043
rect 4893 3003 4951 3009
rect 5350 3000 5356 3052
rect 5408 3040 5414 3052
rect 5813 3043 5871 3049
rect 5813 3040 5825 3043
rect 5408 3012 5825 3040
rect 5408 3000 5414 3012
rect 5813 3009 5825 3012
rect 5859 3009 5871 3043
rect 5813 3003 5871 3009
rect 5902 3000 5908 3052
rect 5960 3040 5966 3052
rect 6365 3043 6423 3049
rect 6365 3040 6377 3043
rect 5960 3012 6377 3040
rect 5960 3000 5966 3012
rect 6365 3009 6377 3012
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 7193 3043 7251 3049
rect 7193 3040 7205 3043
rect 6512 3012 7205 3040
rect 6512 3000 6518 3012
rect 7193 3009 7205 3012
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 7742 3000 7748 3052
rect 7800 3040 7806 3052
rect 8772 3049 8800 3080
rect 9030 3068 9036 3120
rect 9088 3108 9094 3120
rect 9088 3080 10088 3108
rect 9088 3068 9094 3080
rect 8481 3043 8539 3049
rect 8481 3040 8493 3043
rect 7800 3012 8493 3040
rect 7800 3000 7806 3012
rect 8481 3009 8493 3012
rect 8527 3009 8539 3043
rect 8481 3003 8539 3009
rect 8757 3043 8815 3049
rect 8757 3009 8769 3043
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 8846 3000 8852 3052
rect 8904 3040 8910 3052
rect 10060 3049 10088 3080
rect 12158 3068 12164 3120
rect 12216 3108 12222 3120
rect 12216 3080 13308 3108
rect 12216 3068 12222 3080
rect 9677 3043 9735 3049
rect 9677 3040 9689 3043
rect 8904 3012 9689 3040
rect 8904 3000 8910 3012
rect 9677 3009 9689 3012
rect 9723 3009 9735 3043
rect 9677 3003 9735 3009
rect 10045 3043 10103 3049
rect 10045 3009 10057 3043
rect 10091 3009 10103 3043
rect 10045 3003 10103 3009
rect 10686 3000 10692 3052
rect 10744 3040 10750 3052
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 10744 3012 11713 3040
rect 10744 3000 10750 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 11790 3000 11796 3052
rect 11848 3040 11854 3052
rect 13280 3049 13308 3080
rect 13814 3068 13820 3120
rect 13872 3108 13878 3120
rect 15102 3108 15108 3120
rect 13872 3080 15108 3108
rect 13872 3068 13878 3080
rect 15102 3068 15108 3080
rect 15160 3068 15166 3120
rect 12897 3043 12955 3049
rect 12897 3040 12909 3043
rect 11848 3012 12909 3040
rect 11848 3000 11854 3012
rect 12897 3009 12909 3012
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 13265 3043 13323 3049
rect 13265 3009 13277 3043
rect 13311 3009 13323 3043
rect 13265 3003 13323 3009
rect 14182 3000 14188 3052
rect 14240 3040 14246 3052
rect 15764 3049 15792 3148
rect 17310 3136 17316 3188
rect 17368 3176 17374 3188
rect 19058 3176 19064 3188
rect 17368 3148 19064 3176
rect 17368 3136 17374 3148
rect 19058 3136 19064 3148
rect 19116 3136 19122 3188
rect 19702 3136 19708 3188
rect 19760 3176 19766 3188
rect 34330 3176 34336 3188
rect 19760 3148 21496 3176
rect 19760 3136 19766 3148
rect 16206 3068 16212 3120
rect 16264 3108 16270 3120
rect 16264 3080 17724 3108
rect 16264 3068 16270 3080
rect 15381 3043 15439 3049
rect 15381 3040 15393 3043
rect 14240 3012 15393 3040
rect 14240 3000 14246 3012
rect 15381 3009 15393 3012
rect 15427 3009 15439 3043
rect 15381 3003 15439 3009
rect 15749 3043 15807 3049
rect 15749 3009 15761 3043
rect 15795 3009 15807 3043
rect 15749 3003 15807 3009
rect 16022 3000 16028 3052
rect 16080 3040 16086 3052
rect 17696 3049 17724 3080
rect 18598 3068 18604 3120
rect 18656 3108 18662 3120
rect 18656 3080 20208 3108
rect 18656 3068 18662 3080
rect 17405 3043 17463 3049
rect 17405 3040 17417 3043
rect 16080 3012 17417 3040
rect 16080 3000 16086 3012
rect 17405 3009 17417 3012
rect 17451 3009 17463 3043
rect 17405 3003 17463 3009
rect 17681 3043 17739 3049
rect 17681 3009 17693 3043
rect 17727 3009 17739 3043
rect 17681 3003 17739 3009
rect 18046 3000 18052 3052
rect 18104 3040 18110 3052
rect 20180 3049 20208 3080
rect 19521 3043 19579 3049
rect 19521 3040 19533 3043
rect 18104 3012 19533 3040
rect 18104 3000 18110 3012
rect 19521 3009 19533 3012
rect 19567 3009 19579 3043
rect 19521 3003 19579 3009
rect 20165 3043 20223 3049
rect 20165 3009 20177 3043
rect 20211 3009 20223 3043
rect 20165 3003 20223 3009
rect 20254 3000 20260 3052
rect 20312 3040 20318 3052
rect 21468 3049 21496 3148
rect 31864 3148 34336 3176
rect 21634 3068 21640 3120
rect 21692 3108 21698 3120
rect 21692 3080 22968 3108
rect 21692 3068 21698 3080
rect 21085 3043 21143 3049
rect 21085 3040 21097 3043
rect 20312 3012 21097 3040
rect 20312 3000 20318 3012
rect 21085 3009 21097 3012
rect 21131 3009 21143 3043
rect 21085 3003 21143 3009
rect 21453 3043 21511 3049
rect 21453 3009 21465 3043
rect 21499 3009 21511 3043
rect 21453 3003 21511 3009
rect 22097 3043 22155 3049
rect 22097 3009 22109 3043
rect 22143 3040 22155 3043
rect 22186 3040 22192 3052
rect 22143 3012 22192 3040
rect 22143 3009 22155 3012
rect 22097 3003 22155 3009
rect 22186 3000 22192 3012
rect 22244 3000 22250 3052
rect 22554 3000 22560 3052
rect 22612 3040 22618 3052
rect 22940 3049 22968 3080
rect 22649 3043 22707 3049
rect 22649 3040 22661 3043
rect 22612 3012 22661 3040
rect 22612 3000 22618 3012
rect 22649 3009 22661 3012
rect 22695 3009 22707 3043
rect 22649 3003 22707 3009
rect 22925 3043 22983 3049
rect 22925 3009 22937 3043
rect 22971 3009 22983 3043
rect 22925 3003 22983 3009
rect 24305 3043 24363 3049
rect 24305 3009 24317 3043
rect 24351 3040 24363 3043
rect 24486 3040 24492 3052
rect 24351 3012 24492 3040
rect 24351 3009 24363 3012
rect 24305 3003 24363 3009
rect 24486 3000 24492 3012
rect 24544 3000 24550 3052
rect 25593 3043 25651 3049
rect 25593 3009 25605 3043
rect 25639 3040 25651 3043
rect 25774 3040 25780 3052
rect 25639 3012 25780 3040
rect 25639 3009 25651 3012
rect 25593 3003 25651 3009
rect 25774 3000 25780 3012
rect 25832 3000 25838 3052
rect 27982 3000 27988 3052
rect 28040 3040 28046 3052
rect 28169 3043 28227 3049
rect 28169 3040 28181 3043
rect 28040 3012 28181 3040
rect 28040 3000 28046 3012
rect 28169 3009 28181 3012
rect 28215 3009 28227 3043
rect 28169 3003 28227 3009
rect 28445 3043 28503 3049
rect 28445 3009 28457 3043
rect 28491 3040 28503 3043
rect 28718 3040 28724 3052
rect 28491 3012 28724 3040
rect 28491 3009 28503 3012
rect 28445 3003 28503 3009
rect 28718 3000 28724 3012
rect 28776 3000 28782 3052
rect 31570 3040 31576 3052
rect 31531 3012 31576 3040
rect 31570 3000 31576 3012
rect 31628 3000 31634 3052
rect 31864 3049 31892 3148
rect 34330 3136 34336 3148
rect 34388 3136 34394 3188
rect 36630 3176 36636 3188
rect 34532 3148 36636 3176
rect 34422 3108 34428 3120
rect 32876 3080 34428 3108
rect 31849 3043 31907 3049
rect 31849 3009 31861 3043
rect 31895 3009 31907 3043
rect 31849 3003 31907 3009
rect 32401 3043 32459 3049
rect 32401 3009 32413 3043
rect 32447 3040 32459 3043
rect 32766 3040 32772 3052
rect 32447 3012 32772 3040
rect 32447 3009 32459 3012
rect 32401 3003 32459 3009
rect 32766 3000 32772 3012
rect 32824 3000 32830 3052
rect 32876 3049 32904 3080
rect 34422 3068 34428 3080
rect 34480 3068 34486 3120
rect 32861 3043 32919 3049
rect 32861 3009 32873 3043
rect 32907 3009 32919 3043
rect 32861 3003 32919 3009
rect 33137 3043 33195 3049
rect 33137 3009 33149 3043
rect 33183 3040 33195 3043
rect 33226 3040 33232 3052
rect 33183 3012 33232 3040
rect 33183 3009 33195 3012
rect 33137 3003 33195 3009
rect 33226 3000 33232 3012
rect 33284 3000 33290 3052
rect 33689 3043 33747 3049
rect 33689 3009 33701 3043
rect 33735 3040 33747 3043
rect 33778 3040 33784 3052
rect 33735 3012 33784 3040
rect 33735 3009 33747 3012
rect 33689 3003 33747 3009
rect 33778 3000 33784 3012
rect 33836 3000 33842 3052
rect 34532 3049 34560 3148
rect 36630 3136 36636 3148
rect 36688 3136 36694 3188
rect 36817 3179 36875 3185
rect 36817 3145 36829 3179
rect 36863 3176 36875 3179
rect 38470 3176 38476 3188
rect 36863 3148 38476 3176
rect 36863 3145 36875 3148
rect 36817 3139 36875 3145
rect 38470 3136 38476 3148
rect 38528 3136 38534 3188
rect 38654 3136 38660 3188
rect 38712 3176 38718 3188
rect 39574 3176 39580 3188
rect 38712 3148 39580 3176
rect 38712 3136 38718 3148
rect 39574 3136 39580 3148
rect 39632 3136 39638 3188
rect 42150 3176 42156 3188
rect 40420 3148 42156 3176
rect 37734 3108 37740 3120
rect 35728 3080 37740 3108
rect 35728 3049 35756 3080
rect 37734 3068 37740 3080
rect 37792 3068 37798 3120
rect 39022 3108 39028 3120
rect 37844 3080 39028 3108
rect 34517 3043 34575 3049
rect 34517 3009 34529 3043
rect 34563 3009 34575 3043
rect 34517 3003 34575 3009
rect 35713 3043 35771 3049
rect 35713 3009 35725 3043
rect 35759 3009 35771 3043
rect 35713 3003 35771 3009
rect 35989 3043 36047 3049
rect 35989 3009 36001 3043
rect 36035 3040 36047 3043
rect 37550 3040 37556 3052
rect 36035 3012 37556 3040
rect 36035 3009 36047 3012
rect 35989 3003 36047 3009
rect 37550 3000 37556 3012
rect 37608 3000 37614 3052
rect 2406 2932 2412 2984
rect 2464 2972 2470 2984
rect 3053 2975 3111 2981
rect 3053 2972 3065 2975
rect 2464 2944 3065 2972
rect 2464 2932 2470 2944
rect 3053 2941 3065 2944
rect 3099 2941 3111 2975
rect 3053 2935 3111 2941
rect 3234 2932 3240 2984
rect 3292 2972 3298 2984
rect 3329 2975 3387 2981
rect 3329 2972 3341 2975
rect 3292 2944 3341 2972
rect 3292 2932 3298 2944
rect 3329 2941 3341 2944
rect 3375 2941 3387 2975
rect 3329 2935 3387 2941
rect 4798 2932 4804 2984
rect 4856 2972 4862 2984
rect 5169 2975 5227 2981
rect 5169 2972 5181 2975
rect 4856 2944 5181 2972
rect 4856 2932 4862 2944
rect 5169 2941 5181 2944
rect 5215 2941 5227 2975
rect 5169 2935 5227 2941
rect 6086 2932 6092 2984
rect 6144 2972 6150 2984
rect 6641 2975 6699 2981
rect 6641 2972 6653 2975
rect 6144 2944 6653 2972
rect 6144 2932 6150 2944
rect 6641 2941 6653 2944
rect 6687 2941 6699 2975
rect 6641 2935 6699 2941
rect 6914 2932 6920 2984
rect 6972 2972 6978 2984
rect 7469 2975 7527 2981
rect 7469 2972 7481 2975
rect 6972 2944 7481 2972
rect 6972 2932 6978 2944
rect 7469 2941 7481 2944
rect 7515 2941 7527 2975
rect 7469 2935 7527 2941
rect 7558 2932 7564 2984
rect 7616 2972 7622 2984
rect 9033 2975 9091 2981
rect 9033 2972 9045 2975
rect 7616 2944 9045 2972
rect 7616 2932 7622 2944
rect 9033 2941 9045 2944
rect 9079 2941 9091 2975
rect 9033 2935 9091 2941
rect 9398 2932 9404 2984
rect 9456 2972 9462 2984
rect 10321 2975 10379 2981
rect 10321 2972 10333 2975
rect 9456 2944 10333 2972
rect 9456 2932 9462 2944
rect 10321 2941 10333 2944
rect 10367 2941 10379 2975
rect 10321 2935 10379 2941
rect 10410 2932 10416 2984
rect 10468 2972 10474 2984
rect 11333 2975 11391 2981
rect 11333 2972 11345 2975
rect 10468 2944 11345 2972
rect 10468 2932 10474 2944
rect 11333 2941 11345 2944
rect 11379 2941 11391 2975
rect 11333 2935 11391 2941
rect 11514 2932 11520 2984
rect 11572 2972 11578 2984
rect 11572 2944 12480 2972
rect 11572 2932 11578 2944
rect 1949 2907 2007 2913
rect 1949 2873 1961 2907
rect 1995 2904 2007 2907
rect 2774 2904 2780 2916
rect 1995 2876 2780 2904
rect 1995 2873 2007 2876
rect 1949 2867 2007 2873
rect 2774 2864 2780 2876
rect 2832 2864 2838 2916
rect 3510 2904 3516 2916
rect 2976 2876 3516 2904
rect 1118 2796 1124 2848
rect 1176 2836 1182 2848
rect 2225 2839 2283 2845
rect 2225 2836 2237 2839
rect 1176 2808 2237 2836
rect 1176 2796 1182 2808
rect 2225 2805 2237 2808
rect 2271 2805 2283 2839
rect 2225 2799 2283 2805
rect 2501 2839 2559 2845
rect 2501 2805 2513 2839
rect 2547 2836 2559 2839
rect 2976 2836 3004 2876
rect 3510 2864 3516 2876
rect 3568 2864 3574 2916
rect 7190 2864 7196 2916
rect 7248 2904 7254 2916
rect 7929 2907 7987 2913
rect 7929 2904 7941 2907
rect 7248 2876 7941 2904
rect 7248 2864 7254 2876
rect 7929 2873 7941 2876
rect 7975 2873 7987 2907
rect 7929 2867 7987 2873
rect 8478 2864 8484 2916
rect 8536 2904 8542 2916
rect 9309 2907 9367 2913
rect 9309 2904 9321 2907
rect 8536 2876 9321 2904
rect 8536 2864 8542 2876
rect 9309 2873 9321 2876
rect 9355 2873 9367 2907
rect 9309 2867 9367 2873
rect 9674 2864 9680 2916
rect 9732 2904 9738 2916
rect 10597 2907 10655 2913
rect 10597 2904 10609 2907
rect 9732 2876 10609 2904
rect 9732 2864 9738 2876
rect 10597 2873 10609 2876
rect 10643 2873 10655 2907
rect 10597 2867 10655 2873
rect 11238 2864 11244 2916
rect 11296 2904 11302 2916
rect 12253 2907 12311 2913
rect 12253 2904 12265 2907
rect 11296 2876 12265 2904
rect 11296 2864 11302 2876
rect 12253 2873 12265 2876
rect 12299 2873 12311 2907
rect 12253 2867 12311 2873
rect 2547 2808 3004 2836
rect 2547 2805 2559 2808
rect 2501 2799 2559 2805
rect 5166 2796 5172 2848
rect 5224 2836 5230 2848
rect 5537 2839 5595 2845
rect 5537 2836 5549 2839
rect 5224 2808 5549 2836
rect 5224 2796 5230 2808
rect 5537 2805 5549 2808
rect 5583 2805 5595 2839
rect 5537 2799 5595 2805
rect 5626 2796 5632 2848
rect 5684 2836 5690 2848
rect 6089 2839 6147 2845
rect 6089 2836 6101 2839
rect 5684 2808 6101 2836
rect 5684 2796 5690 2808
rect 6089 2805 6101 2808
rect 6135 2805 6147 2839
rect 6089 2799 6147 2805
rect 7006 2796 7012 2848
rect 7064 2836 7070 2848
rect 8205 2839 8263 2845
rect 8205 2836 8217 2839
rect 7064 2808 8217 2836
rect 7064 2796 7070 2808
rect 8205 2805 8217 2808
rect 8251 2805 8263 2839
rect 8205 2799 8263 2805
rect 9950 2796 9956 2848
rect 10008 2836 10014 2848
rect 10965 2839 11023 2845
rect 10965 2836 10977 2839
rect 10008 2808 10977 2836
rect 10008 2796 10014 2808
rect 10965 2805 10977 2808
rect 11011 2805 11023 2839
rect 10965 2799 11023 2805
rect 11054 2796 11060 2848
rect 11112 2836 11118 2848
rect 11977 2839 12035 2845
rect 11977 2836 11989 2839
rect 11112 2808 11989 2836
rect 11112 2796 11118 2808
rect 11977 2805 11989 2808
rect 12023 2805 12035 2839
rect 12452 2836 12480 2944
rect 12526 2932 12532 2984
rect 12584 2972 12590 2984
rect 13633 2975 13691 2981
rect 13633 2972 13645 2975
rect 12584 2944 13645 2972
rect 12584 2932 12590 2944
rect 13633 2941 13645 2944
rect 13679 2941 13691 2975
rect 13633 2935 13691 2941
rect 13814 2932 13820 2984
rect 13872 2972 13878 2984
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 13872 2944 14841 2972
rect 13872 2932 13878 2944
rect 14829 2941 14841 2944
rect 14875 2941 14887 2975
rect 14829 2935 14887 2941
rect 14918 2932 14924 2984
rect 14976 2972 14982 2984
rect 16209 2975 16267 2981
rect 16209 2972 16221 2975
rect 14976 2944 16221 2972
rect 14976 2932 14982 2944
rect 16209 2941 16221 2944
rect 16255 2941 16267 2975
rect 16758 2972 16764 2984
rect 16719 2944 16764 2972
rect 16209 2935 16267 2941
rect 16758 2932 16764 2944
rect 16816 2932 16822 2984
rect 18414 2932 18420 2984
rect 18472 2972 18478 2984
rect 19889 2975 19947 2981
rect 19889 2972 19901 2975
rect 18472 2944 19901 2972
rect 18472 2932 18478 2944
rect 19889 2941 19901 2944
rect 19935 2941 19947 2975
rect 19889 2935 19947 2941
rect 20438 2932 20444 2984
rect 20496 2972 20502 2984
rect 21821 2975 21879 2981
rect 21821 2972 21833 2975
rect 20496 2944 21833 2972
rect 20496 2932 20502 2944
rect 21821 2941 21833 2944
rect 21867 2941 21879 2975
rect 21821 2935 21879 2941
rect 22462 2932 22468 2984
rect 22520 2972 22526 2984
rect 23569 2975 23627 2981
rect 23569 2972 23581 2975
rect 22520 2944 23581 2972
rect 22520 2932 22526 2944
rect 23569 2941 23581 2944
rect 23615 2941 23627 2975
rect 23569 2935 23627 2941
rect 32125 2975 32183 2981
rect 32125 2941 32137 2975
rect 32171 2972 32183 2975
rect 33413 2975 33471 2981
rect 32171 2944 33364 2972
rect 32171 2941 32183 2944
rect 32125 2935 32183 2941
rect 13078 2864 13084 2916
rect 13136 2904 13142 2916
rect 14277 2907 14335 2913
rect 14277 2904 14289 2907
rect 13136 2876 14289 2904
rect 13136 2864 13142 2876
rect 14277 2873 14289 2876
rect 14323 2873 14335 2907
rect 15102 2904 15108 2916
rect 15063 2876 15108 2904
rect 14277 2867 14335 2873
rect 15102 2864 15108 2876
rect 15160 2864 15166 2916
rect 15654 2864 15660 2916
rect 15712 2904 15718 2916
rect 17037 2907 17095 2913
rect 17037 2904 17049 2907
rect 15712 2876 17049 2904
rect 15712 2864 15718 2876
rect 17037 2873 17049 2876
rect 17083 2873 17095 2907
rect 17037 2867 17095 2873
rect 17126 2864 17132 2916
rect 17184 2904 17190 2916
rect 18601 2907 18659 2913
rect 18601 2904 18613 2907
rect 17184 2876 18613 2904
rect 17184 2864 17190 2876
rect 18601 2873 18613 2876
rect 18647 2873 18659 2907
rect 18874 2904 18880 2916
rect 18835 2876 18880 2904
rect 18601 2867 18659 2873
rect 18874 2864 18880 2876
rect 18932 2864 18938 2916
rect 18966 2864 18972 2916
rect 19024 2904 19030 2916
rect 20533 2907 20591 2913
rect 20533 2904 20545 2907
rect 19024 2876 20545 2904
rect 19024 2864 19030 2876
rect 20533 2873 20545 2876
rect 20579 2873 20591 2907
rect 20533 2867 20591 2873
rect 20990 2864 20996 2916
rect 21048 2904 21054 2916
rect 22373 2907 22431 2913
rect 22373 2904 22385 2907
rect 21048 2876 22385 2904
rect 21048 2864 21054 2876
rect 22373 2873 22385 2876
rect 22419 2873 22431 2907
rect 23201 2907 23259 2913
rect 23201 2904 23213 2907
rect 22373 2867 22431 2873
rect 22480 2876 23213 2904
rect 12529 2839 12587 2845
rect 12529 2836 12541 2839
rect 12452 2808 12541 2836
rect 11977 2799 12035 2805
rect 12529 2805 12541 2808
rect 12575 2805 12587 2839
rect 12529 2799 12587 2805
rect 12710 2796 12716 2848
rect 12768 2836 12774 2848
rect 13909 2839 13967 2845
rect 13909 2836 13921 2839
rect 12768 2808 13921 2836
rect 12768 2796 12774 2808
rect 13909 2805 13921 2808
rect 13955 2805 13967 2839
rect 13909 2799 13967 2805
rect 14185 2839 14243 2845
rect 14185 2805 14197 2839
rect 14231 2836 14243 2839
rect 14553 2839 14611 2845
rect 14553 2836 14565 2839
rect 14231 2808 14565 2836
rect 14231 2805 14243 2808
rect 14185 2799 14243 2805
rect 14553 2805 14565 2808
rect 14599 2805 14611 2839
rect 14553 2799 14611 2805
rect 14642 2796 14648 2848
rect 14700 2836 14706 2848
rect 16485 2839 16543 2845
rect 16485 2836 16497 2839
rect 14700 2808 16497 2836
rect 14700 2796 14706 2808
rect 16485 2805 16497 2808
rect 16531 2805 16543 2839
rect 16485 2799 16543 2805
rect 16574 2796 16580 2848
rect 16632 2836 16638 2848
rect 18049 2839 18107 2845
rect 18049 2836 18061 2839
rect 16632 2808 18061 2836
rect 16632 2796 16638 2808
rect 18049 2805 18061 2808
rect 18095 2805 18107 2839
rect 18049 2799 18107 2805
rect 19058 2796 19064 2848
rect 19116 2836 19122 2848
rect 19153 2839 19211 2845
rect 19153 2836 19165 2839
rect 19116 2808 19165 2836
rect 19116 2796 19122 2808
rect 19153 2805 19165 2808
rect 19199 2805 19211 2839
rect 19153 2799 19211 2805
rect 19242 2796 19248 2848
rect 19300 2836 19306 2848
rect 20809 2839 20867 2845
rect 20809 2836 20821 2839
rect 19300 2808 20821 2836
rect 19300 2796 19306 2808
rect 20809 2805 20821 2808
rect 20855 2805 20867 2839
rect 20809 2799 20867 2805
rect 20898 2796 20904 2848
rect 20956 2836 20962 2848
rect 22480 2836 22508 2876
rect 23201 2873 23213 2876
rect 23247 2873 23259 2907
rect 23201 2867 23259 2873
rect 28721 2907 28779 2913
rect 28721 2873 28733 2907
rect 28767 2904 28779 2907
rect 29270 2904 29276 2916
rect 28767 2876 29276 2904
rect 28767 2873 28779 2876
rect 28721 2867 28779 2873
rect 29270 2864 29276 2876
rect 29328 2864 29334 2916
rect 30653 2907 30711 2913
rect 30653 2873 30665 2907
rect 30699 2904 30711 2907
rect 32398 2904 32404 2916
rect 30699 2876 32404 2904
rect 30699 2873 30711 2876
rect 30653 2867 30711 2873
rect 32398 2864 32404 2876
rect 32456 2864 32462 2916
rect 33336 2904 33364 2944
rect 33413 2941 33425 2975
rect 33459 2972 33471 2975
rect 35158 2972 35164 2984
rect 33459 2944 35164 2972
rect 33459 2941 33471 2944
rect 33413 2935 33471 2941
rect 35158 2932 35164 2944
rect 35216 2932 35222 2984
rect 35253 2975 35311 2981
rect 35253 2941 35265 2975
rect 35299 2972 35311 2975
rect 37182 2972 37188 2984
rect 35299 2944 37188 2972
rect 35299 2941 35311 2944
rect 35253 2935 35311 2941
rect 37182 2932 37188 2944
rect 37240 2932 37246 2984
rect 34241 2907 34299 2913
rect 33336 2876 33456 2904
rect 20956 2808 22508 2836
rect 23845 2839 23903 2845
rect 20956 2796 20962 2808
rect 23845 2805 23857 2839
rect 23891 2836 23903 2839
rect 25866 2836 25872 2848
rect 23891 2808 25872 2836
rect 23891 2805 23903 2808
rect 23845 2799 23903 2805
rect 25866 2796 25872 2808
rect 25924 2796 25930 2848
rect 33428 2836 33456 2876
rect 34241 2873 34253 2907
rect 34287 2904 34299 2907
rect 34977 2907 35035 2913
rect 34287 2876 34928 2904
rect 34287 2873 34299 2876
rect 34241 2867 34299 2873
rect 34790 2836 34796 2848
rect 33428 2808 34796 2836
rect 34790 2796 34796 2808
rect 34848 2796 34854 2848
rect 34900 2836 34928 2876
rect 34977 2873 34989 2907
rect 35023 2904 35035 2907
rect 35023 2876 35756 2904
rect 35023 2873 35035 2876
rect 34977 2867 35035 2873
rect 35618 2836 35624 2848
rect 34900 2808 35624 2836
rect 35618 2796 35624 2808
rect 35676 2796 35682 2848
rect 35728 2836 35756 2876
rect 35802 2864 35808 2916
rect 35860 2904 35866 2916
rect 36446 2904 36452 2916
rect 35860 2876 36452 2904
rect 35860 2864 35866 2876
rect 36446 2864 36452 2876
rect 36504 2864 36510 2916
rect 36541 2907 36599 2913
rect 36541 2873 36553 2907
rect 36587 2904 36599 2907
rect 36817 2907 36875 2913
rect 36817 2904 36829 2907
rect 36587 2876 36829 2904
rect 36587 2873 36599 2876
rect 36541 2867 36599 2873
rect 36817 2873 36829 2876
rect 36863 2873 36875 2907
rect 36817 2867 36875 2873
rect 36906 2864 36912 2916
rect 36964 2904 36970 2916
rect 37844 2904 37872 3080
rect 39022 3068 39028 3080
rect 39080 3068 39086 3120
rect 37921 3043 37979 3049
rect 37921 3009 37933 3043
rect 37967 3040 37979 3043
rect 39390 3040 39396 3052
rect 37967 3012 39396 3040
rect 37967 3009 37979 3012
rect 37921 3003 37979 3009
rect 39390 3000 39396 3012
rect 39448 3000 39454 3052
rect 39482 3000 39488 3052
rect 39540 3040 39546 3052
rect 40420 3049 40448 3148
rect 42150 3136 42156 3148
rect 42208 3136 42214 3188
rect 44358 3176 44364 3188
rect 42904 3148 44364 3176
rect 42518 3108 42524 3120
rect 40788 3080 42524 3108
rect 40788 3049 40816 3080
rect 42518 3068 42524 3080
rect 42576 3068 42582 3120
rect 40405 3043 40463 3049
rect 39540 3012 40356 3040
rect 39540 3000 39546 3012
rect 38565 2975 38623 2981
rect 38565 2941 38577 2975
rect 38611 2972 38623 2975
rect 40126 2972 40132 2984
rect 38611 2944 40132 2972
rect 38611 2941 38623 2944
rect 38565 2935 38623 2941
rect 40126 2932 40132 2944
rect 40184 2932 40190 2984
rect 40328 2972 40356 3012
rect 40405 3009 40417 3043
rect 40451 3009 40463 3043
rect 40405 3003 40463 3009
rect 40773 3043 40831 3049
rect 40773 3009 40785 3043
rect 40819 3009 40831 3043
rect 40773 3003 40831 3009
rect 41049 3043 41107 3049
rect 41049 3009 41061 3043
rect 41095 3040 41107 3043
rect 41966 3040 41972 3052
rect 41095 3012 41972 3040
rect 41095 3009 41107 3012
rect 41049 3003 41107 3009
rect 41966 3000 41972 3012
rect 42024 3000 42030 3052
rect 42153 3043 42211 3049
rect 42153 3009 42165 3043
rect 42199 3040 42211 3043
rect 42794 3040 42800 3052
rect 42199 3012 42800 3040
rect 42199 3009 42211 3012
rect 42153 3003 42211 3009
rect 42794 3000 42800 3012
rect 42852 3000 42858 3052
rect 42904 3049 42932 3148
rect 44358 3136 44364 3148
rect 44416 3136 44422 3188
rect 46198 3176 46204 3188
rect 44836 3148 46204 3176
rect 44542 3108 44548 3120
rect 43180 3080 44548 3108
rect 43180 3049 43208 3080
rect 44542 3068 44548 3080
rect 44600 3068 44606 3120
rect 42889 3043 42947 3049
rect 42889 3009 42901 3043
rect 42935 3009 42947 3043
rect 42889 3003 42947 3009
rect 43165 3043 43223 3049
rect 43165 3009 43177 3043
rect 43211 3009 43223 3043
rect 43165 3003 43223 3009
rect 43625 3043 43683 3049
rect 43625 3009 43637 3043
rect 43671 3040 43683 3043
rect 44266 3040 44272 3052
rect 43671 3012 44272 3040
rect 43671 3009 43683 3012
rect 43625 3003 43683 3009
rect 44266 3000 44272 3012
rect 44324 3000 44330 3052
rect 44836 3049 44864 3148
rect 46198 3136 46204 3148
rect 46256 3136 46262 3188
rect 58894 3176 58900 3188
rect 56244 3148 58900 3176
rect 45833 3111 45891 3117
rect 45833 3077 45845 3111
rect 45879 3108 45891 3111
rect 46934 3108 46940 3120
rect 45879 3080 46940 3108
rect 45879 3077 45891 3080
rect 45833 3071 45891 3077
rect 46934 3068 46940 3080
rect 46992 3068 46998 3120
rect 48590 3108 48596 3120
rect 47320 3080 48596 3108
rect 44821 3043 44879 3049
rect 44821 3009 44833 3043
rect 44867 3009 44879 3043
rect 44821 3003 44879 3009
rect 45281 3043 45339 3049
rect 45281 3009 45293 3043
rect 45327 3040 45339 3043
rect 46750 3040 46756 3052
rect 45327 3012 46756 3040
rect 45327 3009 45339 3012
rect 45281 3003 45339 3009
rect 46750 3000 46756 3012
rect 46808 3000 46814 3052
rect 47320 3049 47348 3080
rect 48590 3068 48596 3080
rect 48648 3068 48654 3120
rect 50430 3108 50436 3120
rect 49344 3080 50436 3108
rect 47305 3043 47363 3049
rect 47305 3009 47317 3043
rect 47351 3009 47363 3043
rect 47305 3003 47363 3009
rect 47581 3043 47639 3049
rect 47581 3009 47593 3043
rect 47627 3040 47639 3043
rect 48038 3040 48044 3052
rect 47627 3012 48044 3040
rect 47627 3009 47639 3012
rect 47581 3003 47639 3009
rect 48038 3000 48044 3012
rect 48096 3000 48102 3052
rect 48317 3043 48375 3049
rect 48317 3009 48329 3043
rect 48363 3040 48375 3043
rect 48958 3040 48964 3052
rect 48363 3012 48964 3040
rect 48363 3009 48375 3012
rect 48317 3003 48375 3009
rect 48958 3000 48964 3012
rect 49016 3000 49022 3052
rect 49344 3049 49372 3080
rect 50430 3068 50436 3080
rect 50488 3068 50494 3120
rect 51718 3108 51724 3120
rect 50724 3080 51724 3108
rect 49329 3043 49387 3049
rect 49329 3009 49341 3043
rect 49375 3009 49387 3043
rect 49329 3003 49387 3009
rect 49605 3043 49663 3049
rect 49605 3009 49617 3043
rect 49651 3040 49663 3043
rect 50246 3040 50252 3052
rect 49651 3012 50252 3040
rect 49651 3009 49663 3012
rect 49605 3003 49663 3009
rect 50246 3000 50252 3012
rect 50304 3000 50310 3052
rect 50724 3049 50752 3080
rect 51718 3068 51724 3080
rect 51776 3068 51782 3120
rect 52822 3108 52828 3120
rect 52012 3080 52828 3108
rect 50709 3043 50767 3049
rect 50709 3009 50721 3043
rect 50755 3009 50767 3043
rect 50709 3003 50767 3009
rect 50985 3043 51043 3049
rect 50985 3009 50997 3043
rect 51031 3040 51043 3043
rect 51534 3040 51540 3052
rect 51031 3012 51540 3040
rect 51031 3009 51043 3012
rect 50985 3003 51043 3009
rect 51534 3000 51540 3012
rect 51592 3000 51598 3052
rect 52012 3049 52040 3080
rect 52822 3068 52828 3080
rect 52880 3068 52886 3120
rect 54478 3108 54484 3120
rect 53944 3080 54484 3108
rect 51997 3043 52055 3049
rect 51997 3009 52009 3043
rect 52043 3009 52055 3043
rect 51997 3003 52055 3009
rect 53101 3043 53159 3049
rect 53101 3009 53113 3043
rect 53147 3040 53159 3043
rect 53558 3040 53564 3052
rect 53147 3012 53564 3040
rect 53147 3009 53159 3012
rect 53101 3003 53159 3009
rect 53558 3000 53564 3012
rect 53616 3000 53622 3052
rect 53944 3049 53972 3080
rect 54478 3068 54484 3080
rect 54536 3068 54542 3120
rect 53929 3043 53987 3049
rect 53929 3009 53941 3043
rect 53975 3009 53987 3043
rect 53929 3003 53987 3009
rect 54205 3043 54263 3049
rect 54205 3009 54217 3043
rect 54251 3040 54263 3043
rect 54662 3040 54668 3052
rect 54251 3012 54668 3040
rect 54251 3009 54263 3012
rect 54205 3003 54263 3009
rect 54662 3000 54668 3012
rect 54720 3000 54726 3052
rect 55125 3043 55183 3049
rect 55125 3009 55137 3043
rect 55171 3040 55183 3043
rect 55582 3040 55588 3052
rect 55171 3012 55588 3040
rect 55171 3009 55183 3012
rect 55125 3003 55183 3009
rect 55582 3000 55588 3012
rect 55640 3000 55646 3052
rect 56244 3049 56272 3148
rect 58894 3136 58900 3148
rect 58952 3136 58958 3188
rect 58342 3108 58348 3120
rect 56428 3080 58348 3108
rect 56229 3043 56287 3049
rect 56229 3009 56241 3043
rect 56275 3009 56287 3043
rect 56229 3003 56287 3009
rect 41230 2972 41236 2984
rect 40328 2944 41236 2972
rect 41230 2932 41236 2944
rect 41288 2932 41294 2984
rect 41877 2975 41935 2981
rect 41877 2941 41889 2975
rect 41923 2972 41935 2975
rect 43070 2972 43076 2984
rect 41923 2944 43076 2972
rect 41923 2941 41935 2944
rect 41877 2935 41935 2941
rect 43070 2932 43076 2944
rect 43128 2932 43134 2984
rect 44545 2975 44603 2981
rect 44545 2941 44557 2975
rect 44591 2972 44603 2975
rect 45646 2972 45652 2984
rect 44591 2944 45652 2972
rect 44591 2941 44603 2944
rect 44545 2935 44603 2941
rect 45646 2932 45652 2944
rect 45704 2932 45710 2984
rect 46293 2975 46351 2981
rect 46293 2941 46305 2975
rect 46339 2972 46351 2975
rect 47486 2972 47492 2984
rect 46339 2944 47492 2972
rect 46339 2941 46351 2944
rect 46293 2935 46351 2941
rect 47486 2932 47492 2944
rect 47544 2932 47550 2984
rect 48685 2975 48743 2981
rect 48685 2941 48697 2975
rect 48731 2972 48743 2975
rect 49878 2972 49884 2984
rect 48731 2944 49884 2972
rect 48731 2941 48743 2944
rect 48685 2935 48743 2941
rect 49878 2932 49884 2944
rect 49936 2932 49942 2984
rect 49973 2975 50031 2981
rect 49973 2941 49985 2975
rect 50019 2972 50031 2975
rect 50798 2972 50804 2984
rect 50019 2944 50804 2972
rect 50019 2941 50031 2944
rect 49973 2935 50031 2941
rect 50798 2932 50804 2944
rect 50856 2932 50862 2984
rect 51721 2975 51779 2981
rect 51721 2941 51733 2975
rect 51767 2972 51779 2975
rect 52638 2972 52644 2984
rect 51767 2944 52644 2972
rect 51767 2941 51779 2944
rect 51721 2935 51779 2941
rect 52638 2932 52644 2944
rect 52696 2932 52702 2984
rect 52825 2975 52883 2981
rect 52825 2941 52837 2975
rect 52871 2972 52883 2975
rect 53374 2972 53380 2984
rect 52871 2944 53380 2972
rect 52871 2941 52883 2944
rect 52825 2935 52883 2941
rect 53374 2932 53380 2944
rect 53432 2932 53438 2984
rect 54757 2975 54815 2981
rect 54757 2941 54769 2975
rect 54803 2972 54815 2975
rect 55214 2972 55220 2984
rect 54803 2944 55220 2972
rect 54803 2941 54815 2944
rect 54757 2935 54815 2941
rect 55214 2932 55220 2944
rect 55272 2932 55278 2984
rect 55953 2975 56011 2981
rect 55953 2941 55965 2975
rect 55999 2972 56011 2975
rect 56428 2972 56456 3080
rect 58342 3068 58348 3080
rect 58400 3068 58406 3120
rect 56594 3000 56600 3052
rect 56652 3040 56658 3052
rect 56781 3043 56839 3049
rect 56781 3040 56793 3043
rect 56652 3012 56793 3040
rect 56652 3000 56658 3012
rect 56781 3009 56793 3012
rect 56827 3009 56839 3043
rect 56781 3003 56839 3009
rect 57609 3043 57667 3049
rect 57609 3009 57621 3043
rect 57655 3040 57667 3043
rect 58158 3040 58164 3052
rect 57655 3012 58164 3040
rect 57655 3009 57667 3012
rect 57609 3003 57667 3009
rect 58158 3000 58164 3012
rect 58216 3000 58222 3052
rect 55999 2944 56456 2972
rect 55999 2941 56011 2944
rect 55953 2935 56011 2941
rect 56502 2932 56508 2984
rect 56560 2972 56566 2984
rect 57333 2975 57391 2981
rect 57333 2972 57345 2975
rect 56560 2944 57345 2972
rect 56560 2932 56566 2944
rect 57333 2941 57345 2944
rect 57379 2941 57391 2975
rect 57333 2935 57391 2941
rect 36964 2876 37009 2904
rect 37200 2876 37872 2904
rect 38197 2907 38255 2913
rect 36964 2864 36970 2876
rect 36170 2836 36176 2848
rect 35728 2808 36176 2836
rect 36170 2796 36176 2808
rect 36228 2796 36234 2848
rect 36265 2839 36323 2845
rect 36265 2805 36277 2839
rect 36311 2836 36323 2839
rect 37090 2836 37096 2848
rect 36311 2808 37096 2836
rect 36311 2805 36323 2808
rect 36265 2799 36323 2805
rect 37090 2796 37096 2808
rect 37148 2796 37154 2848
rect 37200 2845 37228 2876
rect 38197 2873 38209 2907
rect 38243 2904 38255 2907
rect 39758 2904 39764 2916
rect 38243 2876 39764 2904
rect 38243 2873 38255 2876
rect 38197 2867 38255 2873
rect 39758 2864 39764 2876
rect 39816 2864 39822 2916
rect 40037 2907 40095 2913
rect 40037 2873 40049 2907
rect 40083 2904 40095 2907
rect 41782 2904 41788 2916
rect 40083 2876 41788 2904
rect 40083 2873 40095 2876
rect 40037 2867 40095 2873
rect 41782 2864 41788 2876
rect 41840 2864 41846 2916
rect 42245 2907 42303 2913
rect 42245 2873 42257 2907
rect 42291 2904 42303 2907
rect 43806 2904 43812 2916
rect 42291 2876 43812 2904
rect 42291 2873 42303 2876
rect 42245 2867 42303 2873
rect 43806 2864 43812 2876
rect 43864 2864 43870 2916
rect 43901 2907 43959 2913
rect 43901 2873 43913 2907
rect 43947 2904 43959 2907
rect 44910 2904 44916 2916
rect 43947 2876 44916 2904
rect 43947 2873 43959 2876
rect 43901 2867 43959 2873
rect 44910 2864 44916 2876
rect 44968 2864 44974 2916
rect 45557 2907 45615 2913
rect 45557 2873 45569 2907
rect 45603 2904 45615 2907
rect 45833 2907 45891 2913
rect 45833 2904 45845 2907
rect 45603 2876 45845 2904
rect 45603 2873 45615 2876
rect 45557 2867 45615 2873
rect 45833 2873 45845 2876
rect 45879 2873 45891 2907
rect 45833 2867 45891 2873
rect 46569 2907 46627 2913
rect 46569 2873 46581 2907
rect 46615 2904 46627 2907
rect 47854 2904 47860 2916
rect 46615 2876 47860 2904
rect 46615 2873 46627 2876
rect 46569 2867 46627 2873
rect 47854 2864 47860 2876
rect 47912 2864 47918 2916
rect 48961 2907 49019 2913
rect 48961 2873 48973 2907
rect 49007 2904 49019 2907
rect 49694 2904 49700 2916
rect 49007 2876 49700 2904
rect 49007 2873 49019 2876
rect 48961 2867 49019 2873
rect 49694 2864 49700 2876
rect 49752 2864 49758 2916
rect 50249 2907 50307 2913
rect 50249 2873 50261 2907
rect 50295 2904 50307 2907
rect 50982 2904 50988 2916
rect 50295 2876 50988 2904
rect 50295 2873 50307 2876
rect 50249 2867 50307 2873
rect 50982 2864 50988 2876
rect 51040 2864 51046 2916
rect 51353 2907 51411 2913
rect 51353 2873 51365 2907
rect 51399 2904 51411 2907
rect 52270 2904 52276 2916
rect 51399 2876 52276 2904
rect 51399 2873 51411 2876
rect 51353 2867 51411 2873
rect 52270 2864 52276 2876
rect 52328 2864 52334 2916
rect 52365 2907 52423 2913
rect 52365 2873 52377 2907
rect 52411 2904 52423 2907
rect 53190 2904 53196 2916
rect 52411 2876 53196 2904
rect 52411 2873 52423 2876
rect 52365 2867 52423 2873
rect 53190 2864 53196 2876
rect 53248 2864 53254 2916
rect 53561 2907 53619 2913
rect 53561 2873 53573 2907
rect 53607 2904 53619 2907
rect 54110 2904 54116 2916
rect 53607 2876 54116 2904
rect 53607 2873 53619 2876
rect 53561 2867 53619 2873
rect 54110 2864 54116 2876
rect 54168 2864 54174 2916
rect 54481 2907 54539 2913
rect 54481 2873 54493 2907
rect 54527 2904 54539 2907
rect 55030 2904 55036 2916
rect 54527 2876 55036 2904
rect 54527 2873 54539 2876
rect 54481 2867 54539 2873
rect 55030 2864 55036 2876
rect 55088 2864 55094 2916
rect 55677 2907 55735 2913
rect 55677 2873 55689 2907
rect 55723 2904 55735 2907
rect 56870 2904 56876 2916
rect 55723 2876 56876 2904
rect 55723 2873 55735 2876
rect 55677 2867 55735 2873
rect 56870 2864 56876 2876
rect 56928 2864 56934 2916
rect 57057 2907 57115 2913
rect 57057 2873 57069 2907
rect 57103 2904 57115 2907
rect 57882 2904 57888 2916
rect 57103 2876 57888 2904
rect 57103 2873 57115 2876
rect 57057 2867 57115 2873
rect 57882 2864 57888 2876
rect 57940 2864 57946 2916
rect 37185 2839 37243 2845
rect 37185 2805 37197 2839
rect 37231 2805 37243 2839
rect 37185 2799 37243 2805
rect 37645 2839 37703 2845
rect 37645 2805 37657 2839
rect 37691 2836 37703 2839
rect 38654 2836 38660 2848
rect 37691 2808 38660 2836
rect 37691 2805 37703 2808
rect 37645 2799 37703 2805
rect 38654 2796 38660 2808
rect 38712 2796 38718 2848
rect 38838 2836 38844 2848
rect 38799 2808 38844 2836
rect 38838 2796 38844 2808
rect 38896 2796 38902 2848
rect 39114 2836 39120 2848
rect 39075 2808 39120 2836
rect 39114 2796 39120 2808
rect 39172 2796 39178 2848
rect 39393 2839 39451 2845
rect 39393 2805 39405 2839
rect 39439 2836 39451 2839
rect 39482 2836 39488 2848
rect 39439 2808 39488 2836
rect 39439 2805 39451 2808
rect 39393 2799 39451 2805
rect 39482 2796 39488 2808
rect 39540 2796 39546 2848
rect 39669 2839 39727 2845
rect 39669 2805 39681 2839
rect 39715 2836 39727 2839
rect 41414 2836 41420 2848
rect 39715 2808 41420 2836
rect 39715 2805 39727 2808
rect 39669 2799 39727 2805
rect 41414 2796 41420 2808
rect 41472 2796 41478 2848
rect 41601 2839 41659 2845
rect 41601 2805 41613 2839
rect 41647 2836 41659 2839
rect 42153 2839 42211 2845
rect 42153 2836 42165 2839
rect 41647 2808 42165 2836
rect 41647 2805 41659 2808
rect 41601 2799 41659 2805
rect 42153 2805 42165 2808
rect 42199 2805 42211 2839
rect 42153 2799 42211 2805
rect 42613 2839 42671 2845
rect 42613 2805 42625 2839
rect 42659 2836 42671 2839
rect 44174 2836 44180 2848
rect 42659 2808 44180 2836
rect 42659 2805 42671 2808
rect 42613 2799 42671 2805
rect 44174 2796 44180 2808
rect 44232 2796 44238 2848
rect 44269 2839 44327 2845
rect 44269 2805 44281 2839
rect 44315 2836 44327 2839
rect 45462 2836 45468 2848
rect 44315 2808 45468 2836
rect 44315 2805 44327 2808
rect 44269 2799 44327 2805
rect 45462 2796 45468 2808
rect 45520 2796 45526 2848
rect 46017 2839 46075 2845
rect 46017 2805 46029 2839
rect 46063 2836 46075 2839
rect 47210 2836 47216 2848
rect 46063 2808 47216 2836
rect 46063 2805 46075 2808
rect 46017 2799 46075 2805
rect 47210 2796 47216 2808
rect 47268 2796 47274 2848
rect 48041 2839 48099 2845
rect 48041 2805 48053 2839
rect 48087 2836 48099 2839
rect 49326 2836 49332 2848
rect 48087 2808 49332 2836
rect 48087 2805 48099 2808
rect 48041 2799 48099 2805
rect 49326 2796 49332 2808
rect 49384 2796 49390 2848
rect 56505 2839 56563 2845
rect 56505 2805 56517 2839
rect 56551 2836 56563 2839
rect 59262 2836 59268 2848
rect 56551 2808 59268 2836
rect 56551 2805 56563 2808
rect 56505 2799 56563 2805
rect 59262 2796 59268 2808
rect 59320 2796 59326 2848
rect 1380 2746 58604 2768
rect 1380 2694 11354 2746
rect 11406 2694 27354 2746
rect 27406 2694 43354 2746
rect 43406 2694 58604 2746
rect 1380 2672 58604 2694
rect 1854 2592 1860 2644
rect 1912 2632 1918 2644
rect 2869 2635 2927 2641
rect 2869 2632 2881 2635
rect 1912 2604 2881 2632
rect 1912 2592 1918 2604
rect 2869 2601 2881 2604
rect 2915 2601 2927 2635
rect 3142 2632 3148 2644
rect 3103 2604 3148 2632
rect 2869 2595 2927 2601
rect 3142 2592 3148 2604
rect 3200 2592 3206 2644
rect 4062 2592 4068 2644
rect 4120 2632 4126 2644
rect 4617 2635 4675 2641
rect 4617 2632 4629 2635
rect 4120 2604 4629 2632
rect 4120 2592 4126 2604
rect 4617 2601 4629 2604
rect 4663 2601 4675 2635
rect 4617 2595 4675 2601
rect 8294 2592 8300 2644
rect 8352 2632 8358 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 8352 2604 9137 2632
rect 8352 2592 8358 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9125 2595 9183 2601
rect 10134 2592 10140 2644
rect 10192 2632 10198 2644
rect 11149 2635 11207 2641
rect 11149 2632 11161 2635
rect 10192 2604 11161 2632
rect 10192 2592 10198 2604
rect 11149 2601 11161 2604
rect 11195 2601 11207 2635
rect 11149 2595 11207 2601
rect 11974 2592 11980 2644
rect 12032 2632 12038 2644
rect 13081 2635 13139 2641
rect 13081 2632 13093 2635
rect 12032 2604 13093 2632
rect 12032 2592 12038 2604
rect 13081 2601 13093 2604
rect 13127 2601 13139 2635
rect 13081 2595 13139 2601
rect 15470 2592 15476 2644
rect 15528 2632 15534 2644
rect 16853 2635 16911 2641
rect 16853 2632 16865 2635
rect 15528 2604 16865 2632
rect 15528 2592 15534 2604
rect 16853 2601 16865 2604
rect 16899 2601 16911 2635
rect 16853 2595 16911 2601
rect 17494 2592 17500 2644
rect 17552 2632 17558 2644
rect 18969 2635 19027 2641
rect 18969 2632 18981 2635
rect 17552 2604 18981 2632
rect 17552 2592 17558 2604
rect 18969 2601 18981 2604
rect 19015 2601 19027 2635
rect 18969 2595 19027 2601
rect 21177 2635 21235 2641
rect 21177 2601 21189 2635
rect 21223 2632 21235 2635
rect 21726 2632 21732 2644
rect 21223 2604 21732 2632
rect 21223 2601 21235 2604
rect 21177 2595 21235 2601
rect 21726 2592 21732 2604
rect 21784 2592 21790 2644
rect 22005 2635 22063 2641
rect 22005 2601 22017 2635
rect 22051 2632 22063 2635
rect 22646 2632 22652 2644
rect 22051 2604 22652 2632
rect 22051 2601 22063 2604
rect 22005 2595 22063 2601
rect 22646 2592 22652 2604
rect 22704 2592 22710 2644
rect 23201 2635 23259 2641
rect 23201 2601 23213 2635
rect 23247 2632 23259 2635
rect 23750 2632 23756 2644
rect 23247 2604 23756 2632
rect 23247 2601 23259 2604
rect 23201 2595 23259 2601
rect 23750 2592 23756 2604
rect 23808 2592 23814 2644
rect 23845 2635 23903 2641
rect 23845 2601 23857 2635
rect 23891 2632 23903 2635
rect 23934 2632 23940 2644
rect 23891 2604 23940 2632
rect 23891 2601 23903 2604
rect 23845 2595 23903 2601
rect 23934 2592 23940 2604
rect 23992 2592 23998 2644
rect 24673 2635 24731 2641
rect 24673 2601 24685 2635
rect 24719 2632 24731 2635
rect 24762 2632 24768 2644
rect 24719 2604 24768 2632
rect 24719 2601 24731 2604
rect 24673 2595 24731 2601
rect 24762 2592 24768 2604
rect 24820 2592 24826 2644
rect 24949 2635 25007 2641
rect 24949 2601 24961 2635
rect 24995 2632 25007 2635
rect 25222 2632 25228 2644
rect 24995 2604 25228 2632
rect 24995 2601 25007 2604
rect 24949 2595 25007 2601
rect 25222 2592 25228 2604
rect 25280 2592 25286 2644
rect 25409 2635 25467 2641
rect 25409 2601 25421 2635
rect 25455 2632 25467 2635
rect 25590 2632 25596 2644
rect 25455 2604 25596 2632
rect 25455 2601 25467 2604
rect 25409 2595 25467 2601
rect 25590 2592 25596 2604
rect 25648 2592 25654 2644
rect 25774 2592 25780 2644
rect 25832 2632 25838 2644
rect 25869 2635 25927 2641
rect 25869 2632 25881 2635
rect 25832 2604 25881 2632
rect 25832 2592 25838 2604
rect 25869 2601 25881 2604
rect 25915 2601 25927 2635
rect 25869 2595 25927 2601
rect 26237 2635 26295 2641
rect 26237 2601 26249 2635
rect 26283 2632 26295 2635
rect 26326 2632 26332 2644
rect 26283 2604 26332 2632
rect 26283 2601 26295 2604
rect 26237 2595 26295 2601
rect 26326 2592 26332 2604
rect 26384 2592 26390 2644
rect 26510 2592 26516 2644
rect 26568 2632 26574 2644
rect 26789 2635 26847 2641
rect 26789 2632 26801 2635
rect 26568 2604 26801 2632
rect 26568 2592 26574 2604
rect 26789 2601 26801 2604
rect 26835 2601 26847 2635
rect 27062 2632 27068 2644
rect 27023 2604 27068 2632
rect 26789 2595 26847 2601
rect 27062 2592 27068 2604
rect 27120 2592 27126 2644
rect 27614 2592 27620 2644
rect 27672 2632 27678 2644
rect 27709 2635 27767 2641
rect 27709 2632 27721 2635
rect 27672 2604 27721 2632
rect 27672 2592 27678 2604
rect 27709 2601 27721 2604
rect 27755 2601 27767 2635
rect 27709 2595 27767 2601
rect 28166 2592 28172 2644
rect 28224 2632 28230 2644
rect 28629 2635 28687 2641
rect 28629 2632 28641 2635
rect 28224 2604 28641 2632
rect 28224 2592 28230 2604
rect 28629 2601 28641 2604
rect 28675 2601 28687 2635
rect 28629 2595 28687 2601
rect 29454 2592 29460 2644
rect 29512 2632 29518 2644
rect 29641 2635 29699 2641
rect 29641 2632 29653 2635
rect 29512 2604 29653 2632
rect 29512 2592 29518 2604
rect 29641 2601 29653 2604
rect 29687 2601 29699 2635
rect 29641 2595 29699 2601
rect 29917 2635 29975 2641
rect 29917 2601 29929 2635
rect 29963 2632 29975 2635
rect 30006 2632 30012 2644
rect 29963 2604 30012 2632
rect 29963 2601 29975 2604
rect 29917 2595 29975 2601
rect 30006 2592 30012 2604
rect 30064 2592 30070 2644
rect 30374 2592 30380 2644
rect 30432 2632 30438 2644
rect 30469 2635 30527 2641
rect 30469 2632 30481 2635
rect 30432 2604 30481 2632
rect 30432 2592 30438 2604
rect 30469 2601 30481 2604
rect 30515 2601 30527 2635
rect 30742 2632 30748 2644
rect 30703 2604 30748 2632
rect 30469 2595 30527 2601
rect 30742 2592 30748 2604
rect 30800 2592 30806 2644
rect 31294 2592 31300 2644
rect 31352 2632 31358 2644
rect 31849 2635 31907 2641
rect 31849 2632 31861 2635
rect 31352 2604 31861 2632
rect 31352 2592 31358 2604
rect 31849 2601 31861 2604
rect 31895 2601 31907 2635
rect 33042 2632 33048 2644
rect 33003 2604 33048 2632
rect 31849 2595 31907 2601
rect 33042 2592 33048 2604
rect 33100 2592 33106 2644
rect 33502 2592 33508 2644
rect 33560 2632 33566 2644
rect 34057 2635 34115 2641
rect 34057 2632 34069 2635
rect 33560 2604 34069 2632
rect 33560 2592 33566 2604
rect 34057 2601 34069 2604
rect 34103 2601 34115 2635
rect 34057 2595 34115 2601
rect 34238 2592 34244 2644
rect 34296 2632 34302 2644
rect 34977 2635 35035 2641
rect 34977 2632 34989 2635
rect 34296 2604 34989 2632
rect 34296 2592 34302 2604
rect 34977 2601 34989 2604
rect 35023 2601 35035 2635
rect 34977 2595 35035 2601
rect 35897 2635 35955 2641
rect 35897 2601 35909 2635
rect 35943 2632 35955 2635
rect 37918 2632 37924 2644
rect 35943 2604 37924 2632
rect 35943 2601 35955 2604
rect 35897 2595 35955 2601
rect 37918 2592 37924 2604
rect 37976 2592 37982 2644
rect 38473 2635 38531 2641
rect 38473 2601 38485 2635
rect 38519 2632 38531 2635
rect 40310 2632 40316 2644
rect 38519 2604 40316 2632
rect 38519 2601 38531 2604
rect 38473 2595 38531 2601
rect 40310 2592 40316 2604
rect 40368 2592 40374 2644
rect 41969 2635 42027 2641
rect 41969 2601 41981 2635
rect 42015 2632 42027 2635
rect 43622 2632 43628 2644
rect 42015 2604 43628 2632
rect 42015 2601 42027 2604
rect 41969 2595 42027 2601
rect 43622 2592 43628 2604
rect 43680 2592 43686 2644
rect 45189 2635 45247 2641
rect 45189 2601 45201 2635
rect 45235 2632 45247 2635
rect 46566 2632 46572 2644
rect 45235 2604 46572 2632
rect 45235 2601 45247 2604
rect 45189 2595 45247 2601
rect 46566 2592 46572 2604
rect 46624 2592 46630 2644
rect 47121 2635 47179 2641
rect 47121 2601 47133 2635
rect 47167 2632 47179 2635
rect 48222 2632 48228 2644
rect 47167 2604 48228 2632
rect 47167 2601 47179 2604
rect 47121 2595 47179 2601
rect 48222 2592 48228 2604
rect 48280 2592 48286 2644
rect 50341 2635 50399 2641
rect 50341 2601 50353 2635
rect 50387 2632 50399 2635
rect 50982 2632 50988 2644
rect 50387 2604 50988 2632
rect 50387 2601 50399 2604
rect 50341 2595 50399 2601
rect 50982 2592 50988 2604
rect 51040 2592 51046 2644
rect 51169 2635 51227 2641
rect 51169 2601 51181 2635
rect 51215 2632 51227 2635
rect 52086 2632 52092 2644
rect 51215 2604 52092 2632
rect 51215 2601 51227 2604
rect 51169 2595 51227 2601
rect 52086 2592 52092 2604
rect 52144 2592 52150 2644
rect 53285 2635 53343 2641
rect 53285 2601 53297 2635
rect 53331 2632 53343 2635
rect 53742 2632 53748 2644
rect 53331 2604 53748 2632
rect 53331 2601 53343 2604
rect 53285 2595 53343 2601
rect 53742 2592 53748 2604
rect 53800 2592 53806 2644
rect 55401 2635 55459 2641
rect 55401 2601 55413 2635
rect 55447 2632 55459 2635
rect 55766 2632 55772 2644
rect 55447 2604 55772 2632
rect 55447 2601 55459 2604
rect 55401 2595 55459 2601
rect 55766 2592 55772 2604
rect 55824 2592 55830 2644
rect 56226 2632 56232 2644
rect 56187 2604 56232 2632
rect 56226 2592 56232 2604
rect 56284 2592 56290 2644
rect 56781 2635 56839 2641
rect 56781 2601 56793 2635
rect 56827 2632 56839 2635
rect 57054 2632 57060 2644
rect 56827 2604 57060 2632
rect 56827 2601 56839 2604
rect 56781 2595 56839 2601
rect 57054 2592 57060 2604
rect 57112 2592 57118 2644
rect 566 2524 572 2576
rect 624 2564 630 2576
rect 3421 2567 3479 2573
rect 3421 2564 3433 2567
rect 624 2536 3433 2564
rect 624 2524 630 2536
rect 3421 2533 3433 2536
rect 3467 2533 3479 2567
rect 3421 2527 3479 2533
rect 3970 2524 3976 2576
rect 4028 2564 4034 2576
rect 4341 2567 4399 2573
rect 4341 2564 4353 2567
rect 4028 2536 4353 2564
rect 4028 2524 4034 2536
rect 4341 2533 4353 2536
rect 4387 2533 4399 2567
rect 4341 2527 4399 2533
rect 17862 2524 17868 2576
rect 17920 2564 17926 2576
rect 19337 2567 19395 2573
rect 19337 2564 19349 2567
rect 17920 2536 19349 2564
rect 17920 2524 17926 2536
rect 19337 2533 19349 2536
rect 19383 2533 19395 2567
rect 19337 2527 19395 2533
rect 20533 2567 20591 2573
rect 20533 2533 20545 2567
rect 20579 2564 20591 2567
rect 21358 2564 21364 2576
rect 20579 2536 21364 2564
rect 20579 2533 20591 2536
rect 20533 2527 20591 2533
rect 21358 2524 21364 2536
rect 21416 2524 21422 2576
rect 21545 2567 21603 2573
rect 21545 2533 21557 2567
rect 21591 2564 21603 2567
rect 22278 2564 22284 2576
rect 21591 2536 22284 2564
rect 21591 2533 21603 2536
rect 21545 2527 21603 2533
rect 22278 2524 22284 2536
rect 22336 2524 22342 2576
rect 22741 2567 22799 2573
rect 22741 2533 22753 2567
rect 22787 2564 22799 2567
rect 23382 2564 23388 2576
rect 22787 2536 23388 2564
rect 22787 2533 22799 2536
rect 22741 2527 22799 2533
rect 23382 2524 23388 2536
rect 23440 2524 23446 2576
rect 23569 2567 23627 2573
rect 23569 2533 23581 2567
rect 23615 2564 23627 2567
rect 24118 2564 24124 2576
rect 23615 2536 24124 2564
rect 23615 2533 23627 2536
rect 23569 2527 23627 2533
rect 24118 2524 24124 2536
rect 24176 2524 24182 2576
rect 26050 2564 26056 2576
rect 24228 2536 26056 2564
rect 3050 2456 3056 2508
rect 3108 2496 3114 2508
rect 4893 2499 4951 2505
rect 4893 2496 4905 2499
rect 3108 2468 4905 2496
rect 3108 2456 3114 2468
rect 4893 2465 4905 2468
rect 4939 2465 4951 2499
rect 4893 2459 4951 2465
rect 22465 2499 22523 2505
rect 22465 2465 22477 2499
rect 22511 2496 22523 2499
rect 23198 2496 23204 2508
rect 22511 2468 23204 2496
rect 22511 2465 22523 2468
rect 22465 2459 22523 2465
rect 23198 2456 23204 2468
rect 23256 2456 23262 2508
rect 750 2388 756 2440
rect 808 2428 814 2440
rect 3697 2431 3755 2437
rect 3697 2428 3709 2431
rect 808 2400 3709 2428
rect 808 2388 814 2400
rect 3697 2397 3709 2400
rect 3743 2397 3755 2431
rect 3697 2391 3755 2397
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 20809 2431 20867 2437
rect 20809 2397 20821 2431
rect 20855 2428 20867 2431
rect 21542 2428 21548 2440
rect 20855 2400 21548 2428
rect 20855 2397 20867 2400
rect 20809 2391 20867 2397
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 3988 2360 4016 2391
rect 21542 2388 21548 2400
rect 21600 2388 21606 2440
rect 22922 2388 22928 2440
rect 22980 2428 22986 2440
rect 24228 2428 24256 2536
rect 26050 2524 26056 2536
rect 26108 2524 26114 2576
rect 26142 2524 26148 2576
rect 26200 2564 26206 2576
rect 26418 2564 26424 2576
rect 26200 2536 26424 2564
rect 26200 2524 26206 2536
rect 26418 2524 26424 2536
rect 26476 2524 26482 2576
rect 26878 2524 26884 2576
rect 26936 2564 26942 2576
rect 27341 2567 27399 2573
rect 27341 2564 27353 2567
rect 26936 2536 27353 2564
rect 26936 2524 26942 2536
rect 27341 2533 27353 2536
rect 27387 2533 27399 2567
rect 27341 2527 27399 2533
rect 27522 2524 27528 2576
rect 27580 2564 27586 2576
rect 27985 2567 28043 2573
rect 27985 2564 27997 2567
rect 27580 2536 27997 2564
rect 27580 2524 27586 2536
rect 27985 2533 27997 2536
rect 28031 2533 28043 2567
rect 27985 2527 28043 2533
rect 28353 2567 28411 2573
rect 28353 2533 28365 2567
rect 28399 2564 28411 2567
rect 28902 2564 28908 2576
rect 28399 2536 28908 2564
rect 28399 2533 28411 2536
rect 28353 2527 28411 2533
rect 28902 2524 28908 2536
rect 28960 2524 28966 2576
rect 29365 2567 29423 2573
rect 29365 2533 29377 2567
rect 29411 2564 29423 2567
rect 29822 2564 29828 2576
rect 29411 2536 29828 2564
rect 29411 2533 29423 2536
rect 29365 2527 29423 2533
rect 29822 2524 29828 2536
rect 29880 2524 29886 2576
rect 30193 2567 30251 2573
rect 30193 2533 30205 2567
rect 30239 2564 30251 2567
rect 30558 2564 30564 2576
rect 30239 2536 30564 2564
rect 30239 2533 30251 2536
rect 30193 2527 30251 2533
rect 30558 2524 30564 2536
rect 30616 2524 30622 2576
rect 31662 2524 31668 2576
rect 31720 2564 31726 2576
rect 32401 2567 32459 2573
rect 32401 2564 32413 2567
rect 31720 2536 32413 2564
rect 31720 2524 31726 2536
rect 32401 2533 32413 2536
rect 32447 2533 32459 2567
rect 32401 2527 32459 2533
rect 32677 2567 32735 2573
rect 32677 2533 32689 2567
rect 32723 2564 32735 2567
rect 32950 2564 32956 2576
rect 32723 2536 32956 2564
rect 32723 2533 32735 2536
rect 32677 2527 32735 2533
rect 32950 2524 32956 2536
rect 33008 2524 33014 2576
rect 33686 2524 33692 2576
rect 33744 2564 33750 2576
rect 34333 2567 34391 2573
rect 34333 2564 34345 2567
rect 33744 2536 34345 2564
rect 33744 2524 33750 2536
rect 34333 2533 34345 2536
rect 34379 2533 34391 2567
rect 34333 2527 34391 2533
rect 40957 2567 41015 2573
rect 40957 2533 40969 2567
rect 41003 2564 41015 2567
rect 42702 2564 42708 2576
rect 41003 2536 42708 2564
rect 41003 2533 41015 2536
rect 40957 2527 41015 2533
rect 42702 2524 42708 2536
rect 42760 2524 42766 2576
rect 44545 2567 44603 2573
rect 44545 2533 44557 2567
rect 44591 2564 44603 2567
rect 46014 2564 46020 2576
rect 44591 2536 46020 2564
rect 44591 2533 44603 2536
rect 44545 2527 44603 2533
rect 46014 2524 46020 2536
rect 46072 2524 46078 2576
rect 47857 2567 47915 2573
rect 47857 2533 47869 2567
rect 47903 2564 47915 2567
rect 49142 2564 49148 2576
rect 47903 2536 49148 2564
rect 47903 2533 47915 2536
rect 47857 2527 47915 2533
rect 49142 2524 49148 2536
rect 49200 2524 49206 2576
rect 54849 2567 54907 2573
rect 54849 2533 54861 2567
rect 54895 2564 54907 2567
rect 55950 2564 55956 2576
rect 54895 2536 55956 2564
rect 54895 2533 54907 2536
rect 54849 2527 54907 2533
rect 55950 2524 55956 2536
rect 56008 2524 56014 2576
rect 56505 2567 56563 2573
rect 56505 2533 56517 2567
rect 56551 2564 56563 2567
rect 57606 2564 57612 2576
rect 56551 2536 57612 2564
rect 56551 2533 56563 2536
rect 56505 2527 56563 2533
rect 57606 2524 57612 2536
rect 57664 2524 57670 2576
rect 24305 2499 24363 2505
rect 24305 2465 24317 2499
rect 24351 2496 24363 2499
rect 24670 2496 24676 2508
rect 24351 2468 24676 2496
rect 24351 2465 24363 2468
rect 24305 2459 24363 2465
rect 24670 2456 24676 2468
rect 24728 2456 24734 2508
rect 24762 2456 24768 2508
rect 24820 2496 24826 2508
rect 26234 2496 26240 2508
rect 24820 2468 26240 2496
rect 24820 2456 24826 2468
rect 26234 2456 26240 2468
rect 26292 2456 26298 2508
rect 28258 2496 28264 2508
rect 26344 2468 28264 2496
rect 25498 2428 25504 2440
rect 22980 2400 24256 2428
rect 24320 2400 25504 2428
rect 22980 2388 22986 2400
rect 1360 2332 4016 2360
rect 1360 2320 1366 2332
rect 23106 2320 23112 2372
rect 23164 2360 23170 2372
rect 24320 2360 24348 2400
rect 25498 2388 25504 2400
rect 25556 2388 25562 2440
rect 25590 2388 25596 2440
rect 25648 2428 25654 2440
rect 26344 2428 26372 2468
rect 28258 2456 28264 2468
rect 28316 2456 28322 2508
rect 32214 2456 32220 2508
rect 32272 2496 32278 2508
rect 33597 2499 33655 2505
rect 33597 2496 33609 2499
rect 32272 2468 33609 2496
rect 32272 2456 32278 2468
rect 33597 2465 33609 2468
rect 33643 2465 33655 2499
rect 33597 2459 33655 2465
rect 34054 2456 34060 2508
rect 34112 2496 34118 2508
rect 34701 2499 34759 2505
rect 34701 2496 34713 2499
rect 34112 2468 34713 2496
rect 34112 2456 34118 2468
rect 34701 2465 34713 2468
rect 34747 2465 34759 2499
rect 34701 2459 34759 2465
rect 55125 2499 55183 2505
rect 55125 2465 55137 2499
rect 55171 2496 55183 2499
rect 55171 2468 56272 2496
rect 55171 2465 55183 2468
rect 55125 2459 55183 2465
rect 25648 2400 26372 2428
rect 25648 2388 25654 2400
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 28905 2431 28963 2437
rect 28905 2428 28917 2431
rect 28408 2400 28917 2428
rect 28408 2388 28414 2400
rect 28905 2397 28917 2400
rect 28951 2397 28963 2431
rect 28905 2391 28963 2397
rect 31846 2388 31852 2440
rect 31904 2428 31910 2440
rect 33321 2431 33379 2437
rect 33321 2428 33333 2431
rect 31904 2400 33333 2428
rect 31904 2388 31910 2400
rect 33321 2397 33333 2400
rect 33367 2397 33379 2431
rect 33321 2391 33379 2397
rect 55677 2431 55735 2437
rect 55677 2397 55689 2431
rect 55723 2397 55735 2431
rect 55677 2391 55735 2397
rect 55953 2431 56011 2437
rect 55953 2397 55965 2431
rect 55999 2428 56011 2431
rect 56042 2428 56048 2440
rect 55999 2400 56048 2428
rect 55999 2397 56011 2400
rect 55953 2391 56011 2397
rect 23164 2332 24348 2360
rect 23164 2320 23170 2332
rect 25038 2320 25044 2372
rect 25096 2360 25102 2372
rect 27798 2360 27804 2372
rect 25096 2332 27804 2360
rect 25096 2320 25102 2332
rect 27798 2320 27804 2332
rect 27856 2320 27862 2372
rect 28442 2320 28448 2372
rect 28500 2360 28506 2372
rect 31294 2360 31300 2372
rect 28500 2332 31300 2360
rect 28500 2320 28506 2332
rect 31294 2320 31300 2332
rect 31352 2320 31358 2372
rect 55692 2360 55720 2391
rect 56042 2388 56048 2400
rect 56100 2388 56106 2440
rect 56244 2428 56272 2468
rect 56318 2456 56324 2508
rect 56376 2496 56382 2508
rect 57057 2499 57115 2505
rect 57057 2496 57069 2499
rect 56376 2468 57069 2496
rect 56376 2456 56382 2468
rect 57057 2465 57069 2468
rect 57103 2465 57115 2499
rect 57057 2459 57115 2465
rect 57422 2428 57428 2440
rect 56244 2400 57428 2428
rect 57422 2388 57428 2400
rect 57480 2388 57486 2440
rect 58710 2360 58716 2372
rect 55692 2332 58716 2360
rect 58710 2320 58716 2332
rect 58768 2320 58774 2372
rect 21082 2252 21088 2304
rect 21140 2292 21146 2304
rect 24946 2292 24952 2304
rect 21140 2264 24952 2292
rect 21140 2252 21146 2264
rect 24946 2252 24952 2264
rect 25004 2252 25010 2304
rect 25314 2252 25320 2304
rect 25372 2292 25378 2304
rect 28534 2292 28540 2304
rect 25372 2264 28540 2292
rect 25372 2252 25378 2264
rect 28534 2252 28540 2264
rect 28592 2252 28598 2304
rect 30374 2252 30380 2304
rect 30432 2292 30438 2304
rect 33134 2292 33140 2304
rect 30432 2264 33140 2292
rect 30432 2252 30438 2264
rect 33134 2252 33140 2264
rect 33192 2252 33198 2304
rect 1380 2202 58604 2224
rect 1380 2150 3354 2202
rect 3406 2150 19354 2202
rect 19406 2150 35354 2202
rect 35406 2150 51354 2202
rect 51406 2150 58604 2202
rect 1380 2128 58604 2150
rect 23842 2048 23848 2100
rect 23900 2088 23906 2100
rect 27062 2088 27068 2100
rect 23900 2060 27068 2088
rect 23900 2048 23906 2060
rect 27062 2048 27068 2060
rect 27120 2048 27126 2100
rect 29454 2088 29460 2100
rect 27632 2060 29460 2088
rect 23290 2020 23296 2032
rect 20824 1992 23296 2020
rect 2038 1912 2044 1964
rect 2096 1952 2102 1964
rect 3694 1952 3700 1964
rect 2096 1924 3556 1952
rect 3655 1924 3700 1952
rect 2096 1912 2102 1924
rect 2590 1844 2596 1896
rect 2648 1884 2654 1896
rect 3421 1887 3479 1893
rect 3421 1884 3433 1887
rect 2648 1856 3433 1884
rect 2648 1844 2654 1856
rect 3421 1853 3433 1856
rect 3467 1853 3479 1887
rect 3528 1884 3556 1924
rect 3694 1912 3700 1924
rect 3752 1912 3758 1964
rect 3970 1952 3976 1964
rect 3931 1924 3976 1952
rect 3970 1912 3976 1924
rect 4028 1912 4034 1964
rect 4154 1912 4160 1964
rect 4212 1952 4218 1964
rect 20824 1961 20852 1992
rect 23290 1980 23296 1992
rect 23348 1980 23354 2032
rect 26142 2020 26148 2032
rect 23400 1992 26148 2020
rect 5353 1955 5411 1961
rect 5353 1952 5365 1955
rect 4212 1924 5365 1952
rect 4212 1912 4218 1924
rect 5353 1921 5365 1924
rect 5399 1921 5411 1955
rect 5353 1915 5411 1921
rect 20809 1955 20867 1961
rect 20809 1921 20821 1955
rect 20855 1921 20867 1955
rect 21082 1952 21088 1964
rect 21043 1924 21088 1952
rect 20809 1915 20867 1921
rect 21082 1912 21088 1924
rect 21140 1912 21146 1964
rect 21361 1955 21419 1961
rect 21361 1921 21373 1955
rect 21407 1952 21419 1955
rect 22002 1952 22008 1964
rect 21407 1924 22008 1952
rect 21407 1921 21419 1924
rect 21361 1915 21419 1921
rect 22002 1912 22008 1924
rect 22060 1912 22066 1964
rect 22189 1955 22247 1961
rect 22189 1921 22201 1955
rect 22235 1952 22247 1955
rect 22830 1952 22836 1964
rect 22235 1924 22836 1952
rect 22235 1921 22247 1924
rect 22189 1915 22247 1921
rect 22830 1912 22836 1924
rect 22888 1912 22894 1964
rect 23106 1952 23112 1964
rect 23067 1924 23112 1952
rect 23106 1912 23112 1924
rect 23164 1912 23170 1964
rect 23400 1961 23428 1992
rect 26142 1980 26148 1992
rect 26200 1980 26206 2032
rect 26326 1980 26332 2032
rect 26384 2020 26390 2032
rect 27632 2020 27660 2060
rect 29454 2048 29460 2060
rect 29512 2048 29518 2100
rect 29546 2048 29552 2100
rect 29604 2088 29610 2100
rect 32398 2088 32404 2100
rect 29604 2060 32404 2088
rect 29604 2048 29610 2060
rect 32398 2048 32404 2060
rect 32456 2048 32462 2100
rect 36262 2088 36268 2100
rect 33888 2060 36268 2088
rect 26384 1992 27660 2020
rect 26384 1980 26390 1992
rect 27706 1980 27712 2032
rect 27764 2020 27770 2032
rect 30650 2020 30656 2032
rect 27764 1992 30656 2020
rect 27764 1980 27770 1992
rect 30650 1980 30656 1992
rect 30708 1980 30714 2032
rect 30926 1980 30932 2032
rect 30984 2020 30990 2032
rect 33686 2020 33692 2032
rect 30984 1992 33692 2020
rect 30984 1980 30990 1992
rect 33686 1980 33692 1992
rect 33744 1980 33750 2032
rect 23385 1955 23443 1961
rect 23385 1921 23397 1955
rect 23431 1921 23443 1955
rect 23385 1915 23443 1921
rect 24029 1955 24087 1961
rect 24029 1921 24041 1955
rect 24075 1952 24087 1955
rect 24762 1952 24768 1964
rect 24075 1924 24768 1952
rect 24075 1921 24087 1924
rect 24029 1915 24087 1921
rect 24762 1912 24768 1924
rect 24820 1912 24826 1964
rect 25038 1952 25044 1964
rect 24999 1924 25044 1952
rect 25038 1912 25044 1924
rect 25096 1912 25102 1964
rect 25314 1952 25320 1964
rect 25275 1924 25320 1952
rect 25314 1912 25320 1924
rect 25372 1912 25378 1964
rect 25590 1952 25596 1964
rect 25551 1924 25596 1952
rect 25590 1912 25596 1924
rect 25648 1912 25654 1964
rect 26602 1912 26608 1964
rect 26660 1952 26666 1964
rect 29638 1952 29644 1964
rect 26660 1924 29644 1952
rect 26660 1912 26666 1924
rect 29638 1912 29644 1924
rect 29696 1912 29702 1964
rect 30374 1952 30380 1964
rect 30335 1924 30380 1952
rect 30374 1912 30380 1924
rect 30432 1912 30438 1964
rect 31110 1952 31116 1964
rect 31071 1924 31116 1952
rect 31110 1912 31116 1924
rect 31168 1912 31174 1964
rect 31386 1912 31392 1964
rect 31444 1952 31450 1964
rect 33318 1952 33324 1964
rect 31444 1924 33324 1952
rect 31444 1912 31450 1924
rect 33318 1912 33324 1924
rect 33376 1912 33382 1964
rect 33888 1961 33916 2060
rect 36262 2048 36268 2060
rect 36320 2048 36326 2100
rect 57974 2088 57980 2100
rect 55508 2060 57980 2088
rect 34146 1980 34152 2032
rect 34204 2020 34210 2032
rect 36630 2020 36636 2032
rect 34204 1992 36636 2020
rect 34204 1980 34210 1992
rect 36630 1980 36636 1992
rect 36688 1980 36694 2032
rect 38194 1980 38200 2032
rect 38252 2020 38258 2032
rect 40126 2020 40132 2032
rect 38252 1992 40132 2020
rect 38252 1980 38258 1992
rect 40126 1980 40132 1992
rect 40184 1980 40190 2032
rect 33873 1955 33931 1961
rect 33873 1921 33885 1955
rect 33919 1921 33931 1955
rect 33873 1915 33931 1921
rect 34790 1912 34796 1964
rect 34848 1952 34854 1964
rect 37182 1952 37188 1964
rect 34848 1924 37188 1952
rect 34848 1912 34854 1924
rect 37182 1912 37188 1924
rect 37240 1912 37246 1964
rect 39485 1955 39543 1961
rect 39485 1921 39497 1955
rect 39531 1952 39543 1955
rect 41414 1952 41420 1964
rect 39531 1924 41420 1952
rect 39531 1921 39543 1924
rect 39485 1915 39543 1921
rect 41414 1912 41420 1924
rect 41472 1912 41478 1964
rect 42058 1912 42064 1964
rect 42116 1952 42122 1964
rect 42702 1952 42708 1964
rect 42116 1924 42708 1952
rect 42116 1912 42122 1924
rect 42702 1912 42708 1924
rect 42760 1912 42766 1964
rect 54481 1955 54539 1961
rect 54481 1921 54493 1955
rect 54527 1952 54539 1955
rect 55508 1952 55536 2060
rect 57974 2048 57980 2060
rect 58032 2048 58038 2100
rect 55858 1980 55864 2032
rect 55916 2020 55922 2032
rect 58526 2020 58532 2032
rect 55916 1992 58532 2020
rect 55916 1980 55922 1992
rect 58526 1980 58532 1992
rect 58584 1980 58590 2032
rect 55674 1952 55680 1964
rect 54527 1924 55536 1952
rect 55635 1924 55680 1952
rect 54527 1921 54539 1924
rect 54481 1915 54539 1921
rect 55674 1912 55680 1924
rect 55732 1912 55738 1964
rect 55950 1952 55956 1964
rect 55911 1924 55956 1952
rect 55950 1912 55956 1924
rect 56008 1912 56014 1964
rect 56226 1952 56232 1964
rect 56187 1924 56232 1952
rect 56226 1912 56232 1924
rect 56284 1912 56290 1964
rect 3528 1856 4200 1884
rect 3421 1847 3479 1853
rect 2774 1776 2780 1828
rect 2832 1816 2838 1828
rect 3145 1819 3203 1825
rect 3145 1816 3157 1819
rect 2832 1788 3157 1816
rect 2832 1776 2838 1788
rect 3145 1785 3157 1788
rect 3191 1785 3203 1819
rect 4172 1816 4200 1856
rect 4246 1844 4252 1896
rect 4304 1884 4310 1896
rect 4525 1887 4583 1893
rect 4525 1884 4537 1887
rect 4304 1856 4537 1884
rect 4304 1844 4310 1856
rect 4525 1853 4537 1856
rect 4571 1853 4583 1887
rect 5074 1884 5080 1896
rect 5035 1856 5080 1884
rect 4525 1847 4583 1853
rect 5074 1844 5080 1856
rect 5132 1844 5138 1896
rect 10318 1844 10324 1896
rect 10376 1884 10382 1896
rect 11333 1887 11391 1893
rect 11333 1884 11345 1887
rect 10376 1856 11345 1884
rect 10376 1844 10382 1856
rect 11333 1853 11345 1856
rect 11379 1853 11391 1887
rect 11333 1847 11391 1853
rect 12710 1844 12716 1896
rect 12768 1884 12774 1896
rect 12989 1887 13047 1893
rect 12989 1884 13001 1887
rect 12768 1856 13001 1884
rect 12768 1844 12774 1856
rect 12989 1853 13001 1856
rect 13035 1853 13047 1887
rect 12989 1847 13047 1853
rect 13262 1844 13268 1896
rect 13320 1884 13326 1896
rect 13541 1887 13599 1893
rect 13541 1884 13553 1887
rect 13320 1856 13553 1884
rect 13320 1844 13326 1856
rect 13541 1853 13553 1856
rect 13587 1853 13599 1887
rect 13541 1847 13599 1853
rect 20622 1844 20628 1896
rect 20680 1884 20686 1896
rect 21637 1887 21695 1893
rect 21637 1884 21649 1887
rect 20680 1856 21649 1884
rect 20680 1844 20686 1856
rect 21637 1853 21649 1856
rect 21683 1853 21695 1887
rect 24305 1887 24363 1893
rect 24305 1884 24317 1887
rect 21637 1847 21695 1853
rect 22848 1856 24317 1884
rect 22848 1828 22876 1856
rect 24305 1853 24317 1856
rect 24351 1853 24363 1887
rect 24305 1847 24363 1853
rect 24394 1844 24400 1896
rect 24452 1884 24458 1896
rect 26145 1887 26203 1893
rect 26145 1884 26157 1887
rect 24452 1856 26157 1884
rect 24452 1844 24458 1856
rect 26145 1853 26157 1856
rect 26191 1853 26203 1887
rect 26145 1847 26203 1853
rect 26421 1887 26479 1893
rect 26421 1853 26433 1887
rect 26467 1884 26479 1887
rect 30834 1884 30840 1896
rect 26467 1856 28672 1884
rect 26467 1853 26479 1856
rect 26421 1847 26479 1853
rect 4801 1819 4859 1825
rect 4801 1816 4813 1819
rect 4172 1788 4813 1816
rect 3145 1779 3203 1785
rect 4801 1785 4813 1788
rect 4847 1785 4859 1819
rect 4801 1779 4859 1785
rect 5166 1776 5172 1828
rect 5224 1816 5230 1828
rect 5629 1819 5687 1825
rect 5629 1816 5641 1819
rect 5224 1788 5641 1816
rect 5224 1776 5230 1788
rect 5629 1785 5641 1788
rect 5675 1785 5687 1819
rect 5629 1779 5687 1785
rect 11054 1776 11060 1828
rect 11112 1816 11118 1828
rect 12069 1819 12127 1825
rect 12069 1816 12081 1819
rect 11112 1788 12081 1816
rect 11112 1776 11118 1788
rect 12069 1785 12081 1788
rect 12115 1785 12127 1819
rect 12069 1779 12127 1785
rect 21174 1776 21180 1828
rect 21232 1816 21238 1828
rect 21913 1819 21971 1825
rect 21913 1816 21925 1819
rect 21232 1788 21925 1816
rect 21232 1776 21238 1788
rect 21913 1785 21925 1788
rect 21959 1785 21971 1819
rect 21913 1779 21971 1785
rect 22002 1776 22008 1828
rect 22060 1816 22066 1828
rect 22465 1819 22523 1825
rect 22465 1816 22477 1819
rect 22060 1788 22477 1816
rect 22060 1776 22066 1788
rect 22465 1785 22477 1788
rect 22511 1785 22523 1819
rect 22465 1779 22523 1785
rect 22830 1776 22836 1828
rect 22888 1776 22894 1828
rect 23566 1776 23572 1828
rect 23624 1816 23630 1828
rect 24765 1819 24823 1825
rect 24765 1816 24777 1819
rect 23624 1788 24777 1816
rect 23624 1776 23630 1788
rect 24765 1785 24777 1788
rect 24811 1785 24823 1819
rect 24765 1779 24823 1785
rect 26234 1776 26240 1828
rect 26292 1816 26298 1828
rect 27246 1816 27252 1828
rect 26292 1788 27252 1816
rect 26292 1776 26298 1788
rect 27246 1776 27252 1788
rect 27304 1776 27310 1828
rect 28644 1816 28672 1856
rect 30668 1856 30840 1884
rect 28810 1816 28816 1828
rect 28644 1788 28816 1816
rect 28810 1776 28816 1788
rect 28868 1776 28874 1828
rect 30668 1816 30696 1856
rect 30834 1844 30840 1856
rect 30892 1844 30898 1896
rect 31570 1844 31576 1896
rect 31628 1884 31634 1896
rect 34238 1884 34244 1896
rect 31628 1856 34244 1884
rect 31628 1844 31634 1856
rect 34238 1844 34244 1856
rect 34296 1844 34302 1896
rect 34422 1844 34428 1896
rect 34480 1884 34486 1896
rect 36814 1884 36820 1896
rect 34480 1856 36820 1884
rect 34480 1844 34486 1856
rect 36814 1844 36820 1856
rect 36872 1844 36878 1896
rect 37274 1844 37280 1896
rect 37332 1884 37338 1896
rect 39022 1884 39028 1896
rect 37332 1856 39028 1884
rect 37332 1844 37338 1856
rect 39022 1844 39028 1856
rect 39080 1844 39086 1896
rect 39666 1844 39672 1896
rect 39724 1884 39730 1896
rect 41598 1884 41604 1896
rect 39724 1856 41604 1884
rect 39724 1844 39730 1856
rect 41598 1844 41604 1856
rect 41656 1844 41662 1896
rect 42337 1887 42395 1893
rect 42337 1853 42349 1887
rect 42383 1884 42395 1887
rect 43990 1884 43996 1896
rect 42383 1856 43996 1884
rect 42383 1853 42395 1856
rect 42337 1847 42395 1853
rect 43990 1844 43996 1856
rect 44048 1844 44054 1896
rect 54757 1887 54815 1893
rect 54757 1853 54769 1887
rect 54803 1884 54815 1887
rect 55214 1884 55220 1896
rect 54803 1856 55220 1884
rect 54803 1853 54815 1856
rect 54757 1847 54815 1853
rect 55214 1844 55220 1856
rect 55272 1844 55278 1896
rect 57057 1887 57115 1893
rect 57057 1884 57069 1887
rect 55968 1856 57069 1884
rect 55968 1828 55996 1856
rect 57057 1853 57069 1856
rect 57103 1853 57115 1887
rect 57057 1847 57115 1853
rect 29012 1788 30696 1816
rect 2866 1748 2872 1760
rect 2827 1720 2872 1748
rect 2866 1708 2872 1720
rect 2924 1708 2930 1760
rect 3234 1708 3240 1760
rect 3292 1748 3298 1760
rect 4249 1751 4307 1757
rect 4249 1748 4261 1751
rect 3292 1720 4261 1748
rect 3292 1708 3298 1720
rect 4249 1717 4261 1720
rect 4295 1717 4307 1751
rect 4249 1711 4307 1717
rect 7190 1708 7196 1760
rect 7248 1748 7254 1760
rect 8021 1751 8079 1757
rect 8021 1748 8033 1751
rect 7248 1720 8033 1748
rect 7248 1708 7254 1720
rect 8021 1717 8033 1720
rect 8067 1717 8079 1751
rect 8021 1711 8079 1717
rect 9582 1708 9588 1760
rect 9640 1748 9646 1760
rect 10597 1751 10655 1757
rect 10597 1748 10609 1751
rect 9640 1720 10609 1748
rect 9640 1708 9646 1720
rect 10597 1717 10609 1720
rect 10643 1717 10655 1751
rect 10597 1711 10655 1717
rect 11606 1708 11612 1760
rect 11664 1748 11670 1760
rect 12713 1751 12771 1757
rect 12713 1748 12725 1751
rect 11664 1720 12725 1748
rect 11664 1708 11670 1720
rect 12713 1717 12725 1720
rect 12759 1717 12771 1751
rect 12713 1711 12771 1717
rect 13265 1751 13323 1757
rect 13265 1717 13277 1751
rect 13311 1748 13323 1751
rect 13446 1748 13452 1760
rect 13311 1720 13452 1748
rect 13311 1717 13323 1720
rect 13265 1711 13323 1717
rect 13446 1708 13452 1720
rect 13504 1708 13510 1760
rect 13814 1748 13820 1760
rect 13775 1720 13820 1748
rect 13814 1708 13820 1720
rect 13872 1708 13878 1760
rect 14461 1751 14519 1757
rect 14461 1717 14473 1751
rect 14507 1748 14519 1751
rect 14550 1748 14556 1760
rect 14507 1720 14556 1748
rect 14507 1717 14519 1720
rect 14461 1711 14519 1717
rect 14550 1708 14556 1720
rect 14608 1708 14614 1760
rect 16942 1708 16948 1760
rect 17000 1748 17006 1760
rect 17037 1751 17095 1757
rect 17037 1748 17049 1751
rect 17000 1720 17049 1748
rect 17000 1708 17006 1720
rect 17037 1717 17049 1720
rect 17083 1717 17095 1751
rect 17037 1711 17095 1717
rect 18230 1708 18236 1760
rect 18288 1748 18294 1760
rect 18601 1751 18659 1757
rect 18601 1748 18613 1751
rect 18288 1720 18613 1748
rect 18288 1708 18294 1720
rect 18601 1717 18613 1720
rect 18647 1717 18659 1751
rect 18601 1711 18659 1717
rect 19518 1708 19524 1760
rect 19576 1748 19582 1760
rect 20346 1748 20352 1760
rect 19576 1720 20352 1748
rect 19576 1708 19582 1720
rect 20346 1708 20352 1720
rect 20404 1708 20410 1760
rect 21726 1708 21732 1760
rect 21784 1748 21790 1760
rect 22741 1751 22799 1757
rect 22741 1748 22753 1751
rect 21784 1720 22753 1748
rect 21784 1708 21790 1720
rect 22741 1717 22753 1720
rect 22787 1717 22799 1751
rect 22741 1711 22799 1717
rect 24302 1708 24308 1760
rect 24360 1748 24366 1760
rect 25869 1751 25927 1757
rect 25869 1748 25881 1751
rect 24360 1720 25881 1748
rect 24360 1708 24366 1720
rect 25869 1717 25881 1720
rect 25915 1717 25927 1751
rect 25869 1711 25927 1717
rect 25958 1708 25964 1760
rect 26016 1748 26022 1760
rect 27890 1748 27896 1760
rect 26016 1720 27896 1748
rect 26016 1708 26022 1720
rect 27890 1708 27896 1720
rect 27948 1708 27954 1760
rect 27985 1751 28043 1757
rect 27985 1717 27997 1751
rect 28031 1748 28043 1751
rect 29012 1748 29040 1788
rect 30742 1776 30748 1828
rect 30800 1816 30806 1828
rect 31478 1816 31484 1828
rect 30800 1788 31484 1816
rect 30800 1776 30806 1788
rect 31478 1776 31484 1788
rect 31536 1776 31542 1828
rect 31754 1776 31760 1828
rect 31812 1816 31818 1828
rect 31812 1788 32168 1816
rect 31812 1776 31818 1788
rect 28031 1720 29040 1748
rect 28031 1717 28043 1720
rect 27985 1711 28043 1717
rect 29086 1708 29092 1760
rect 29144 1748 29150 1760
rect 30006 1748 30012 1760
rect 29144 1720 30012 1748
rect 29144 1708 29150 1720
rect 30006 1708 30012 1720
rect 30064 1708 30070 1760
rect 30558 1708 30564 1760
rect 30616 1748 30622 1760
rect 32030 1748 32036 1760
rect 30616 1720 32036 1748
rect 30616 1708 30622 1720
rect 32030 1708 32036 1720
rect 32088 1708 32094 1760
rect 32140 1748 32168 1788
rect 32214 1776 32220 1828
rect 32272 1816 32278 1828
rect 34698 1816 34704 1828
rect 32272 1788 34704 1816
rect 32272 1776 32278 1788
rect 34698 1776 34704 1788
rect 34756 1776 34762 1828
rect 35066 1776 35072 1828
rect 35124 1816 35130 1828
rect 37366 1816 37372 1828
rect 35124 1788 37372 1816
rect 35124 1776 35130 1788
rect 37366 1776 37372 1788
rect 37424 1776 37430 1828
rect 37642 1776 37648 1828
rect 37700 1816 37706 1828
rect 39758 1816 39764 1828
rect 37700 1788 39764 1816
rect 37700 1776 37706 1788
rect 39758 1776 39764 1788
rect 39816 1776 39822 1828
rect 40218 1776 40224 1828
rect 40276 1816 40282 1828
rect 42150 1816 42156 1828
rect 40276 1788 42156 1816
rect 40276 1776 40282 1788
rect 42150 1776 42156 1788
rect 42208 1776 42214 1828
rect 42886 1776 42892 1828
rect 42944 1816 42950 1828
rect 43806 1816 43812 1828
rect 42944 1788 43812 1816
rect 42944 1776 42950 1788
rect 43806 1776 43812 1788
rect 43864 1776 43870 1828
rect 45189 1819 45247 1825
rect 45189 1785 45201 1819
rect 45235 1816 45247 1819
rect 46566 1816 46572 1828
rect 45235 1788 46572 1816
rect 45235 1785 45247 1788
rect 45189 1779 45247 1785
rect 46566 1776 46572 1788
rect 46624 1776 46630 1828
rect 55950 1776 55956 1828
rect 56008 1776 56014 1828
rect 56778 1816 56784 1828
rect 56739 1788 56784 1816
rect 56778 1776 56784 1788
rect 56836 1776 56842 1828
rect 58894 1816 58900 1828
rect 57532 1788 58900 1816
rect 32766 1748 32772 1760
rect 32140 1720 32772 1748
rect 32766 1708 32772 1720
rect 32824 1708 32830 1760
rect 32858 1708 32864 1760
rect 32916 1748 32922 1760
rect 35158 1748 35164 1760
rect 32916 1720 35164 1748
rect 32916 1708 32922 1720
rect 35158 1708 35164 1720
rect 35216 1708 35222 1760
rect 35710 1708 35716 1760
rect 35768 1748 35774 1760
rect 37826 1748 37832 1760
rect 35768 1720 37832 1748
rect 35768 1708 35774 1720
rect 37826 1708 37832 1720
rect 37884 1708 37890 1760
rect 37921 1751 37979 1757
rect 37921 1717 37933 1751
rect 37967 1748 37979 1751
rect 39942 1748 39948 1760
rect 37967 1720 39948 1748
rect 37967 1717 37979 1720
rect 37921 1711 37979 1717
rect 39942 1708 39948 1720
rect 40000 1708 40006 1760
rect 41141 1751 41199 1757
rect 41141 1717 41153 1751
rect 41187 1748 41199 1751
rect 42794 1748 42800 1760
rect 41187 1720 42800 1748
rect 41187 1717 41199 1720
rect 41141 1711 41199 1717
rect 42794 1708 42800 1720
rect 42852 1708 42858 1760
rect 43165 1751 43223 1757
rect 43165 1717 43177 1751
rect 43211 1748 43223 1751
rect 44726 1748 44732 1760
rect 43211 1720 44732 1748
rect 43211 1717 43223 1720
rect 43165 1711 43223 1717
rect 44726 1708 44732 1720
rect 44784 1708 44790 1760
rect 45462 1708 45468 1760
rect 45520 1748 45526 1760
rect 46934 1748 46940 1760
rect 45520 1720 46940 1748
rect 45520 1708 45526 1720
rect 46934 1708 46940 1720
rect 46992 1708 46998 1760
rect 48317 1751 48375 1757
rect 48317 1717 48329 1751
rect 48363 1748 48375 1751
rect 49510 1748 49516 1760
rect 48363 1720 49516 1748
rect 48363 1717 48375 1720
rect 48317 1711 48375 1717
rect 49510 1708 49516 1720
rect 49568 1708 49574 1760
rect 49973 1751 50031 1757
rect 49973 1717 49985 1751
rect 50019 1748 50031 1751
rect 50982 1748 50988 1760
rect 50019 1720 50988 1748
rect 50019 1717 50031 1720
rect 49973 1711 50031 1717
rect 50982 1708 50988 1720
rect 51040 1708 51046 1760
rect 55217 1751 55275 1757
rect 55217 1717 55229 1751
rect 55263 1748 55275 1751
rect 55582 1748 55588 1760
rect 55263 1720 55588 1748
rect 55263 1717 55275 1720
rect 55217 1711 55275 1717
rect 55582 1708 55588 1720
rect 55640 1708 55646 1760
rect 56502 1748 56508 1760
rect 56463 1720 56508 1748
rect 56502 1708 56508 1720
rect 56560 1708 56566 1760
rect 56594 1708 56600 1760
rect 56652 1748 56658 1760
rect 57532 1748 57560 1788
rect 58894 1776 58900 1788
rect 58952 1776 58958 1828
rect 56652 1720 57560 1748
rect 57609 1751 57667 1757
rect 56652 1708 56658 1720
rect 57609 1717 57621 1751
rect 57655 1748 57667 1751
rect 59078 1748 59084 1760
rect 57655 1720 59084 1748
rect 57655 1717 57667 1720
rect 57609 1711 57667 1717
rect 59078 1708 59084 1720
rect 59136 1708 59142 1760
rect 1380 1658 58604 1680
rect 1380 1606 11354 1658
rect 11406 1606 27354 1658
rect 27406 1606 43354 1658
rect 43406 1606 58604 1658
rect 1380 1584 58604 1606
rect 566 1504 572 1556
rect 624 1544 630 1556
rect 2869 1547 2927 1553
rect 2869 1544 2881 1547
rect 624 1516 2881 1544
rect 624 1504 630 1516
rect 2869 1513 2881 1516
rect 2915 1513 2927 1547
rect 2869 1507 2927 1513
rect 3878 1504 3884 1556
rect 3936 1544 3942 1556
rect 4617 1547 4675 1553
rect 4617 1544 4629 1547
rect 3936 1516 4629 1544
rect 3936 1504 3942 1516
rect 4617 1513 4629 1516
rect 4663 1513 4675 1547
rect 4617 1507 4675 1513
rect 6638 1504 6644 1556
rect 6696 1544 6702 1556
rect 7837 1547 7895 1553
rect 7837 1544 7849 1547
rect 6696 1516 7849 1544
rect 6696 1504 6702 1516
rect 7837 1513 7849 1516
rect 7883 1513 7895 1547
rect 7837 1507 7895 1513
rect 8110 1504 8116 1556
rect 8168 1544 8174 1556
rect 8168 1516 8340 1544
rect 8168 1504 8174 1516
rect 1486 1436 1492 1488
rect 1544 1476 1550 1488
rect 2041 1479 2099 1485
rect 2041 1476 2053 1479
rect 1544 1448 2053 1476
rect 1544 1436 1550 1448
rect 2041 1445 2053 1448
rect 2087 1445 2099 1479
rect 3421 1479 3479 1485
rect 3421 1476 3433 1479
rect 2041 1439 2099 1445
rect 2700 1448 3433 1476
rect 1302 1368 1308 1420
rect 1360 1408 1366 1420
rect 1360 1380 1808 1408
rect 1360 1368 1366 1380
rect 1780 1340 1808 1380
rect 1854 1368 1860 1420
rect 1912 1408 1918 1420
rect 2317 1411 2375 1417
rect 2317 1408 2329 1411
rect 1912 1380 2329 1408
rect 1912 1368 1918 1380
rect 2317 1377 2329 1380
rect 2363 1377 2375 1411
rect 2317 1371 2375 1377
rect 2406 1368 2412 1420
rect 2464 1408 2470 1420
rect 2593 1411 2651 1417
rect 2593 1408 2605 1411
rect 2464 1380 2605 1408
rect 2464 1368 2470 1380
rect 2593 1377 2605 1380
rect 2639 1377 2651 1411
rect 2593 1371 2651 1377
rect 2700 1340 2728 1448
rect 3421 1445 3433 1448
rect 3467 1445 3479 1479
rect 3421 1439 3479 1445
rect 3694 1436 3700 1488
rect 3752 1476 3758 1488
rect 3973 1479 4031 1485
rect 3973 1476 3985 1479
rect 3752 1448 3985 1476
rect 3752 1436 3758 1448
rect 3973 1445 3985 1448
rect 4019 1445 4031 1479
rect 3973 1439 4031 1445
rect 4798 1436 4804 1488
rect 4856 1476 4862 1488
rect 5629 1479 5687 1485
rect 5629 1476 5641 1479
rect 4856 1448 5641 1476
rect 4856 1436 4862 1448
rect 5629 1445 5641 1448
rect 5675 1445 5687 1479
rect 5629 1439 5687 1445
rect 5718 1436 5724 1488
rect 5776 1476 5782 1488
rect 6273 1479 6331 1485
rect 6273 1476 6285 1479
rect 5776 1448 6285 1476
rect 5776 1436 5782 1448
rect 6273 1445 6285 1448
rect 6319 1445 6331 1479
rect 6273 1439 6331 1445
rect 6362 1436 6368 1488
rect 6420 1476 6426 1488
rect 7193 1479 7251 1485
rect 7193 1476 7205 1479
rect 6420 1448 7205 1476
rect 6420 1436 6426 1448
rect 7193 1445 7205 1448
rect 7239 1445 7251 1479
rect 7193 1439 7251 1445
rect 7374 1436 7380 1488
rect 7432 1476 7438 1488
rect 8205 1479 8263 1485
rect 8205 1476 8217 1479
rect 7432 1448 8217 1476
rect 7432 1436 7438 1448
rect 8205 1445 8217 1448
rect 8251 1445 8263 1479
rect 8312 1476 8340 1516
rect 8478 1504 8484 1556
rect 8536 1544 8542 1556
rect 9309 1547 9367 1553
rect 9309 1544 9321 1547
rect 8536 1516 9321 1544
rect 8536 1504 8542 1516
rect 9309 1513 9321 1516
rect 9355 1513 9367 1547
rect 9309 1507 9367 1513
rect 9766 1504 9772 1556
rect 9824 1544 9830 1556
rect 11241 1547 11299 1553
rect 11241 1544 11253 1547
rect 9824 1516 11253 1544
rect 9824 1504 9830 1516
rect 11241 1513 11253 1516
rect 11287 1513 11299 1547
rect 11241 1507 11299 1513
rect 11514 1504 11520 1556
rect 11572 1544 11578 1556
rect 12345 1547 12403 1553
rect 12345 1544 12357 1547
rect 11572 1516 12357 1544
rect 11572 1504 11578 1516
rect 12345 1513 12357 1516
rect 12391 1513 12403 1547
rect 12345 1507 12403 1513
rect 12621 1547 12679 1553
rect 12621 1513 12633 1547
rect 12667 1544 12679 1547
rect 13449 1547 13507 1553
rect 13449 1544 13461 1547
rect 12667 1516 13461 1544
rect 12667 1513 12679 1516
rect 12621 1507 12679 1513
rect 13449 1513 13461 1516
rect 13495 1513 13507 1547
rect 13449 1507 13507 1513
rect 13998 1504 14004 1556
rect 14056 1544 14062 1556
rect 14277 1547 14335 1553
rect 14277 1544 14289 1547
rect 14056 1516 14289 1544
rect 14056 1504 14062 1516
rect 14277 1513 14289 1516
rect 14323 1513 14335 1547
rect 14277 1507 14335 1513
rect 18782 1504 18788 1556
rect 18840 1544 18846 1556
rect 19705 1547 19763 1553
rect 19705 1544 19717 1547
rect 18840 1516 19717 1544
rect 18840 1504 18846 1516
rect 19705 1513 19717 1516
rect 19751 1513 19763 1547
rect 19705 1507 19763 1513
rect 20070 1504 20076 1556
rect 20128 1544 20134 1556
rect 20901 1547 20959 1553
rect 20901 1544 20913 1547
rect 20128 1516 20913 1544
rect 20128 1504 20134 1516
rect 20901 1513 20913 1516
rect 20947 1513 20959 1547
rect 22922 1544 22928 1556
rect 22883 1516 22928 1544
rect 20901 1507 20959 1513
rect 22922 1504 22928 1516
rect 22980 1504 22986 1556
rect 23014 1504 23020 1556
rect 23072 1544 23078 1556
rect 24305 1547 24363 1553
rect 24305 1544 24317 1547
rect 23072 1516 24317 1544
rect 23072 1504 23078 1516
rect 24305 1513 24317 1516
rect 24351 1513 24363 1547
rect 24305 1507 24363 1513
rect 24857 1547 24915 1553
rect 24857 1513 24869 1547
rect 24903 1544 24915 1547
rect 25038 1544 25044 1556
rect 24903 1516 25044 1544
rect 24903 1513 24915 1516
rect 24857 1507 24915 1513
rect 25038 1504 25044 1516
rect 25096 1504 25102 1556
rect 25133 1547 25191 1553
rect 25133 1513 25145 1547
rect 25179 1544 25191 1547
rect 27614 1544 27620 1556
rect 25179 1516 27620 1544
rect 25179 1513 25191 1516
rect 25133 1507 25191 1513
rect 27614 1504 27620 1516
rect 27672 1504 27678 1556
rect 27706 1504 27712 1556
rect 27764 1544 27770 1556
rect 28353 1547 28411 1553
rect 27764 1516 27809 1544
rect 27764 1504 27770 1516
rect 28353 1513 28365 1547
rect 28399 1544 28411 1547
rect 28442 1544 28448 1556
rect 28399 1516 28448 1544
rect 28399 1513 28411 1516
rect 28353 1507 28411 1513
rect 28442 1504 28448 1516
rect 28500 1504 28506 1556
rect 29086 1544 29092 1556
rect 28552 1516 29092 1544
rect 9033 1479 9091 1485
rect 9033 1476 9045 1479
rect 8312 1448 9045 1476
rect 8205 1439 8263 1445
rect 9033 1445 9045 1448
rect 9079 1445 9091 1479
rect 9033 1439 9091 1445
rect 9214 1436 9220 1488
rect 9272 1476 9278 1488
rect 10229 1479 10287 1485
rect 10229 1476 10241 1479
rect 9272 1448 10241 1476
rect 9272 1436 9278 1448
rect 10229 1445 10241 1448
rect 10275 1445 10287 1479
rect 10229 1439 10287 1445
rect 10870 1436 10876 1488
rect 10928 1476 10934 1488
rect 11885 1479 11943 1485
rect 11885 1476 11897 1479
rect 10928 1448 11897 1476
rect 10928 1436 10934 1448
rect 11885 1445 11897 1448
rect 11931 1445 11943 1479
rect 11885 1439 11943 1445
rect 12158 1436 12164 1488
rect 12216 1476 12222 1488
rect 13173 1479 13231 1485
rect 13173 1476 13185 1479
rect 12216 1448 13185 1476
rect 12216 1436 12222 1448
rect 13173 1445 13185 1448
rect 13219 1445 13231 1479
rect 13173 1439 13231 1445
rect 16206 1436 16212 1488
rect 16264 1476 16270 1488
rect 16945 1479 17003 1485
rect 16945 1476 16957 1479
rect 16264 1448 16957 1476
rect 16264 1436 16270 1448
rect 16945 1445 16957 1448
rect 16991 1445 17003 1479
rect 16945 1439 17003 1445
rect 17678 1436 17684 1488
rect 17736 1476 17742 1488
rect 18049 1479 18107 1485
rect 18049 1476 18061 1479
rect 17736 1448 18061 1476
rect 17736 1436 17742 1448
rect 18049 1445 18061 1448
rect 18095 1445 18107 1479
rect 18049 1439 18107 1445
rect 18598 1436 18604 1488
rect 18656 1476 18662 1488
rect 19061 1479 19119 1485
rect 19061 1476 19073 1479
rect 18656 1448 19073 1476
rect 18656 1436 18662 1448
rect 19061 1445 19073 1448
rect 19107 1445 19119 1479
rect 19061 1439 19119 1445
rect 19886 1436 19892 1488
rect 19944 1476 19950 1488
rect 20625 1479 20683 1485
rect 20625 1476 20637 1479
rect 19944 1448 20637 1476
rect 19944 1436 19950 1448
rect 20625 1445 20637 1448
rect 20671 1445 20683 1479
rect 21453 1479 21511 1485
rect 21453 1476 21465 1479
rect 20625 1439 20683 1445
rect 20732 1448 21465 1476
rect 3145 1411 3203 1417
rect 3145 1377 3157 1411
rect 3191 1408 3203 1411
rect 3234 1408 3240 1420
rect 3191 1380 3240 1408
rect 3191 1377 3203 1380
rect 3145 1371 3203 1377
rect 3234 1368 3240 1380
rect 3292 1368 3298 1420
rect 3510 1368 3516 1420
rect 3568 1408 3574 1420
rect 4341 1411 4399 1417
rect 4341 1408 4353 1411
rect 3568 1380 3740 1408
rect 3568 1368 3574 1380
rect 3712 1349 3740 1380
rect 3804 1380 4353 1408
rect 1780 1312 2728 1340
rect 3697 1343 3755 1349
rect 3697 1309 3709 1343
rect 3743 1309 3755 1343
rect 3697 1303 3755 1309
rect 934 1232 940 1284
rect 992 1272 998 1284
rect 3804 1272 3832 1380
rect 4341 1377 4353 1380
rect 4387 1377 4399 1411
rect 4341 1371 4399 1377
rect 4430 1368 4436 1420
rect 4488 1408 4494 1420
rect 4893 1411 4951 1417
rect 4893 1408 4905 1411
rect 4488 1380 4905 1408
rect 4488 1368 4494 1380
rect 4893 1377 4905 1380
rect 4939 1377 4951 1411
rect 4893 1371 4951 1377
rect 4982 1368 4988 1420
rect 5040 1408 5046 1420
rect 5353 1411 5411 1417
rect 5353 1408 5365 1411
rect 5040 1380 5365 1408
rect 5040 1368 5046 1380
rect 5353 1377 5365 1380
rect 5399 1377 5411 1411
rect 5353 1371 5411 1377
rect 5534 1368 5540 1420
rect 5592 1408 5598 1420
rect 5997 1411 6055 1417
rect 5997 1408 6009 1411
rect 5592 1380 6009 1408
rect 5592 1368 5598 1380
rect 5997 1377 6009 1380
rect 6043 1377 6055 1411
rect 5997 1371 6055 1377
rect 6086 1368 6092 1420
rect 6144 1408 6150 1420
rect 6641 1411 6699 1417
rect 6641 1408 6653 1411
rect 6144 1380 6653 1408
rect 6144 1368 6150 1380
rect 6641 1377 6653 1380
rect 6687 1377 6699 1411
rect 6641 1371 6699 1377
rect 6822 1368 6828 1420
rect 6880 1408 6886 1420
rect 7561 1411 7619 1417
rect 7561 1408 7573 1411
rect 6880 1380 7573 1408
rect 6880 1368 6886 1380
rect 7561 1377 7573 1380
rect 7607 1377 7619 1411
rect 7561 1371 7619 1377
rect 7926 1368 7932 1420
rect 7984 1408 7990 1420
rect 8757 1411 8815 1417
rect 8757 1408 8769 1411
rect 7984 1380 8769 1408
rect 7984 1368 7990 1380
rect 8757 1377 8769 1380
rect 8803 1377 8815 1411
rect 8757 1371 8815 1377
rect 8846 1368 8852 1420
rect 8904 1408 8910 1420
rect 9585 1411 9643 1417
rect 9585 1408 9597 1411
rect 8904 1380 9597 1408
rect 8904 1368 8910 1380
rect 9585 1377 9597 1380
rect 9631 1377 9643 1411
rect 9585 1371 9643 1377
rect 9950 1368 9956 1420
rect 10008 1408 10014 1420
rect 10965 1411 11023 1417
rect 10965 1408 10977 1411
rect 10008 1380 10977 1408
rect 10008 1368 10014 1380
rect 10965 1377 10977 1380
rect 11011 1377 11023 1411
rect 11517 1411 11575 1417
rect 11517 1408 11529 1411
rect 10965 1371 11023 1377
rect 11072 1380 11529 1408
rect 7650 1300 7656 1352
rect 7708 1340 7714 1352
rect 8481 1343 8539 1349
rect 8481 1340 8493 1343
rect 7708 1312 8493 1340
rect 7708 1300 7714 1312
rect 8481 1309 8493 1312
rect 8527 1309 8539 1343
rect 8481 1303 8539 1309
rect 9030 1300 9036 1352
rect 9088 1340 9094 1352
rect 10505 1343 10563 1349
rect 10505 1340 10517 1343
rect 9088 1312 10517 1340
rect 9088 1300 9094 1312
rect 10505 1309 10517 1312
rect 10551 1309 10563 1343
rect 10505 1303 10563 1309
rect 10594 1300 10600 1352
rect 10652 1340 10658 1352
rect 11072 1340 11100 1380
rect 11517 1377 11529 1380
rect 11563 1377 11575 1411
rect 11517 1371 11575 1377
rect 11974 1368 11980 1420
rect 12032 1408 12038 1420
rect 12032 1380 12296 1408
rect 12032 1368 12038 1380
rect 10652 1312 11100 1340
rect 12268 1340 12296 1380
rect 12342 1368 12348 1420
rect 12400 1408 12406 1420
rect 12621 1411 12679 1417
rect 12621 1408 12633 1411
rect 12400 1380 12633 1408
rect 12400 1368 12406 1380
rect 12621 1377 12633 1380
rect 12667 1377 12679 1411
rect 12894 1408 12900 1420
rect 12855 1380 12900 1408
rect 12621 1371 12679 1377
rect 12894 1368 12900 1380
rect 12952 1368 12958 1420
rect 13725 1411 13783 1417
rect 13725 1408 13737 1411
rect 13004 1380 13737 1408
rect 13004 1340 13032 1380
rect 13725 1377 13737 1380
rect 13771 1377 13783 1411
rect 13725 1371 13783 1377
rect 14001 1411 14059 1417
rect 14001 1377 14013 1411
rect 14047 1408 14059 1411
rect 14182 1408 14188 1420
rect 14047 1380 14188 1408
rect 14047 1377 14059 1380
rect 14001 1371 14059 1377
rect 14182 1368 14188 1380
rect 14240 1368 14246 1420
rect 14645 1411 14703 1417
rect 14645 1377 14657 1411
rect 14691 1408 14703 1411
rect 14734 1408 14740 1420
rect 14691 1380 14740 1408
rect 14691 1377 14703 1380
rect 14645 1371 14703 1377
rect 14734 1368 14740 1380
rect 14792 1368 14798 1420
rect 15013 1411 15071 1417
rect 15013 1377 15025 1411
rect 15059 1408 15071 1411
rect 15102 1408 15108 1420
rect 15059 1380 15108 1408
rect 15059 1377 15071 1380
rect 15013 1371 15071 1377
rect 15102 1368 15108 1380
rect 15160 1368 15166 1420
rect 15286 1408 15292 1420
rect 15247 1380 15292 1408
rect 15286 1368 15292 1380
rect 15344 1368 15350 1420
rect 15654 1368 15660 1420
rect 15712 1408 15718 1420
rect 15749 1411 15807 1417
rect 15749 1408 15761 1411
rect 15712 1380 15761 1408
rect 15712 1368 15718 1380
rect 15749 1377 15761 1380
rect 15795 1377 15807 1411
rect 15749 1371 15807 1377
rect 15838 1368 15844 1420
rect 15896 1408 15902 1420
rect 16025 1411 16083 1417
rect 16025 1408 16037 1411
rect 15896 1380 16037 1408
rect 15896 1368 15902 1380
rect 16025 1377 16037 1380
rect 16071 1377 16083 1411
rect 16390 1408 16396 1420
rect 16351 1380 16396 1408
rect 16025 1371 16083 1377
rect 16390 1368 16396 1380
rect 16448 1368 16454 1420
rect 16574 1368 16580 1420
rect 16632 1408 16638 1420
rect 16669 1411 16727 1417
rect 16669 1408 16681 1411
rect 16632 1380 16681 1408
rect 16632 1368 16638 1380
rect 16669 1377 16681 1380
rect 16715 1377 16727 1411
rect 16669 1371 16727 1377
rect 17126 1368 17132 1420
rect 17184 1408 17190 1420
rect 17313 1411 17371 1417
rect 17313 1408 17325 1411
rect 17184 1380 17325 1408
rect 17184 1368 17190 1380
rect 17313 1377 17325 1380
rect 17359 1377 17371 1411
rect 17313 1371 17371 1377
rect 17494 1368 17500 1420
rect 17552 1408 17558 1420
rect 17773 1411 17831 1417
rect 17773 1408 17785 1411
rect 17552 1380 17785 1408
rect 17552 1368 17558 1380
rect 17773 1377 17785 1380
rect 17819 1377 17831 1411
rect 17773 1371 17831 1377
rect 18138 1368 18144 1420
rect 18196 1408 18202 1420
rect 18196 1380 18644 1408
rect 18196 1368 18202 1380
rect 18616 1349 18644 1380
rect 18966 1368 18972 1420
rect 19024 1408 19030 1420
rect 19429 1411 19487 1417
rect 19429 1408 19441 1411
rect 19024 1380 19441 1408
rect 19024 1368 19030 1380
rect 19429 1377 19441 1380
rect 19475 1377 19487 1411
rect 19429 1371 19487 1377
rect 19518 1368 19524 1420
rect 19576 1408 19582 1420
rect 20073 1411 20131 1417
rect 20073 1408 20085 1411
rect 19576 1380 20085 1408
rect 19576 1368 19582 1380
rect 20073 1377 20085 1380
rect 20119 1377 20131 1411
rect 20346 1408 20352 1420
rect 20307 1380 20352 1408
rect 20073 1371 20131 1377
rect 20346 1368 20352 1380
rect 20404 1368 20410 1420
rect 20438 1368 20444 1420
rect 20496 1408 20502 1420
rect 20732 1408 20760 1448
rect 21453 1445 21465 1448
rect 21499 1445 21511 1479
rect 21453 1439 21511 1445
rect 22278 1436 22284 1488
rect 22336 1476 22342 1488
rect 23385 1479 23443 1485
rect 23385 1476 23397 1479
rect 22336 1448 23397 1476
rect 22336 1436 22342 1448
rect 23385 1445 23397 1448
rect 23431 1445 23443 1479
rect 23385 1439 23443 1445
rect 23750 1436 23756 1488
rect 23808 1476 23814 1488
rect 23808 1448 24716 1476
rect 23808 1436 23814 1448
rect 20496 1380 20760 1408
rect 20496 1368 20502 1380
rect 20990 1368 20996 1420
rect 21048 1408 21054 1420
rect 21913 1411 21971 1417
rect 21913 1408 21925 1411
rect 21048 1380 21925 1408
rect 21048 1368 21054 1380
rect 21913 1377 21925 1380
rect 21959 1377 21971 1411
rect 21913 1371 21971 1377
rect 22557 1411 22615 1417
rect 22557 1377 22569 1411
rect 22603 1408 22615 1411
rect 24581 1411 24639 1417
rect 24581 1408 24593 1411
rect 22603 1380 23336 1408
rect 22603 1377 22615 1380
rect 22557 1371 22615 1377
rect 12268 1312 13032 1340
rect 18601 1343 18659 1349
rect 10652 1300 10658 1312
rect 18601 1309 18613 1343
rect 18647 1309 18659 1343
rect 18601 1303 18659 1309
rect 22281 1343 22339 1349
rect 22281 1309 22293 1343
rect 22327 1309 22339 1343
rect 22281 1303 22339 1309
rect 992 1244 3832 1272
rect 992 1232 998 1244
rect 22296 1204 22324 1303
rect 23308 1272 23336 1380
rect 23400 1380 24593 1408
rect 23400 1352 23428 1380
rect 24581 1377 24593 1380
rect 24627 1377 24639 1411
rect 24688 1408 24716 1448
rect 24762 1436 24768 1488
rect 24820 1476 24826 1488
rect 26053 1479 26111 1485
rect 26053 1476 26065 1479
rect 24820 1448 26065 1476
rect 24820 1436 24826 1448
rect 26053 1445 26065 1448
rect 26099 1445 26111 1479
rect 26326 1476 26332 1488
rect 26287 1448 26332 1476
rect 26053 1439 26111 1445
rect 26326 1436 26332 1448
rect 26384 1436 26390 1488
rect 26602 1476 26608 1488
rect 26563 1448 26608 1476
rect 26602 1436 26608 1448
rect 26660 1436 26666 1488
rect 27157 1479 27215 1485
rect 27157 1445 27169 1479
rect 27203 1476 27215 1479
rect 28552 1476 28580 1516
rect 29086 1504 29092 1516
rect 29144 1504 29150 1556
rect 29181 1547 29239 1553
rect 29181 1513 29193 1547
rect 29227 1544 29239 1547
rect 30558 1544 30564 1556
rect 29227 1516 30564 1544
rect 29227 1513 29239 1516
rect 29181 1507 29239 1513
rect 30558 1504 30564 1516
rect 30616 1504 30622 1556
rect 30653 1547 30711 1553
rect 30653 1513 30665 1547
rect 30699 1544 30711 1547
rect 31386 1544 31392 1556
rect 30699 1516 31392 1544
rect 30699 1513 30711 1516
rect 30653 1507 30711 1513
rect 31386 1504 31392 1516
rect 31444 1504 31450 1556
rect 31570 1544 31576 1556
rect 31531 1516 31576 1544
rect 31570 1504 31576 1516
rect 31628 1504 31634 1556
rect 32214 1544 32220 1556
rect 32175 1516 32220 1544
rect 32214 1504 32220 1516
rect 32272 1504 32278 1556
rect 33778 1544 33784 1556
rect 32416 1516 33784 1544
rect 27203 1448 28580 1476
rect 28629 1479 28687 1485
rect 27203 1445 27215 1448
rect 27157 1439 27215 1445
rect 28629 1445 28641 1479
rect 28675 1476 28687 1479
rect 30742 1476 30748 1488
rect 28675 1448 30748 1476
rect 28675 1445 28687 1448
rect 28629 1439 28687 1445
rect 30742 1436 30748 1448
rect 30800 1436 30806 1488
rect 30926 1476 30932 1488
rect 30887 1448 30932 1476
rect 30926 1436 30932 1448
rect 30984 1436 30990 1488
rect 31205 1479 31263 1485
rect 31205 1445 31217 1479
rect 31251 1476 31263 1479
rect 32416 1476 32444 1516
rect 33778 1504 33784 1516
rect 33836 1504 33842 1556
rect 34146 1544 34152 1556
rect 34107 1516 34152 1544
rect 34146 1504 34152 1516
rect 34204 1504 34210 1556
rect 34422 1544 34428 1556
rect 34383 1516 34428 1544
rect 34422 1504 34428 1516
rect 34480 1504 34486 1556
rect 34790 1544 34796 1556
rect 34751 1516 34796 1544
rect 34790 1504 34796 1516
rect 34848 1504 34854 1556
rect 35066 1544 35072 1556
rect 35027 1516 35072 1544
rect 35066 1504 35072 1516
rect 35124 1504 35130 1556
rect 35526 1544 35532 1556
rect 35268 1516 35532 1544
rect 31251 1448 32444 1476
rect 32493 1479 32551 1485
rect 31251 1445 31263 1448
rect 31205 1439 31263 1445
rect 32493 1445 32505 1479
rect 32539 1476 32551 1479
rect 33873 1479 33931 1485
rect 32539 1448 33548 1476
rect 32539 1445 32551 1448
rect 32493 1439 32551 1445
rect 25409 1411 25467 1417
rect 25409 1408 25421 1411
rect 24688 1380 25421 1408
rect 24581 1371 24639 1377
rect 25409 1377 25421 1380
rect 25455 1377 25467 1411
rect 25409 1371 25467 1377
rect 25777 1411 25835 1417
rect 25777 1377 25789 1411
rect 25823 1408 25835 1411
rect 27985 1411 28043 1417
rect 25823 1380 27936 1408
rect 25823 1377 25835 1380
rect 25777 1371 25835 1377
rect 23382 1300 23388 1352
rect 23440 1300 23446 1352
rect 23753 1343 23811 1349
rect 23753 1309 23765 1343
rect 23799 1340 23811 1343
rect 23842 1340 23848 1352
rect 23799 1312 23848 1340
rect 23799 1309 23811 1312
rect 23753 1303 23811 1309
rect 23842 1300 23848 1312
rect 23900 1300 23906 1352
rect 27433 1343 27491 1349
rect 27433 1309 27445 1343
rect 27479 1309 27491 1343
rect 27433 1303 27491 1309
rect 25774 1272 25780 1284
rect 23308 1244 25780 1272
rect 25774 1232 25780 1244
rect 25832 1232 25838 1284
rect 25406 1204 25412 1216
rect 22296 1176 25412 1204
rect 25406 1164 25412 1176
rect 25464 1164 25470 1216
rect 26142 1164 26148 1216
rect 26200 1204 26206 1216
rect 26694 1204 26700 1216
rect 26200 1176 26700 1204
rect 26200 1164 26206 1176
rect 26694 1164 26700 1176
rect 26752 1164 26758 1216
rect 27448 1204 27476 1303
rect 27908 1272 27936 1380
rect 27985 1377 27997 1411
rect 28031 1408 28043 1411
rect 30190 1408 30196 1420
rect 28031 1380 30196 1408
rect 28031 1377 28043 1380
rect 27985 1371 28043 1377
rect 30190 1368 30196 1380
rect 30248 1368 30254 1420
rect 30285 1411 30343 1417
rect 30285 1377 30297 1411
rect 30331 1408 30343 1411
rect 32582 1408 32588 1420
rect 30331 1380 32588 1408
rect 30331 1377 30343 1380
rect 30285 1371 30343 1377
rect 32582 1368 32588 1380
rect 32640 1368 32646 1420
rect 32858 1408 32864 1420
rect 32819 1380 32864 1408
rect 32858 1368 32864 1380
rect 32916 1368 32922 1420
rect 33229 1411 33287 1417
rect 33229 1377 33241 1411
rect 33275 1408 33287 1411
rect 33275 1380 33456 1408
rect 33275 1377 33287 1380
rect 33229 1371 33287 1377
rect 28905 1343 28963 1349
rect 28905 1309 28917 1343
rect 28951 1309 28963 1343
rect 29546 1340 29552 1352
rect 29507 1312 29552 1340
rect 28905 1303 28963 1309
rect 28810 1272 28816 1284
rect 27908 1244 28816 1272
rect 28810 1232 28816 1244
rect 28868 1232 28874 1284
rect 28920 1272 28948 1303
rect 29546 1300 29552 1312
rect 29604 1300 29610 1352
rect 30009 1343 30067 1349
rect 30009 1309 30021 1343
rect 30055 1340 30067 1343
rect 31754 1340 31760 1352
rect 30055 1312 31760 1340
rect 30055 1309 30067 1312
rect 30009 1303 30067 1309
rect 31754 1300 31760 1312
rect 31812 1300 31818 1352
rect 31849 1343 31907 1349
rect 31849 1309 31861 1343
rect 31895 1309 31907 1343
rect 31849 1303 31907 1309
rect 28920 1244 31800 1272
rect 31772 1216 31800 1244
rect 30374 1204 30380 1216
rect 27448 1176 30380 1204
rect 30374 1164 30380 1176
rect 30432 1164 30438 1216
rect 31754 1164 31760 1216
rect 31812 1164 31818 1216
rect 31864 1204 31892 1303
rect 33428 1272 33456 1380
rect 33520 1340 33548 1448
rect 33873 1445 33885 1479
rect 33919 1476 33931 1479
rect 35268 1476 35296 1516
rect 35526 1504 35532 1516
rect 35584 1504 35590 1556
rect 35710 1544 35716 1556
rect 35671 1516 35716 1544
rect 35710 1504 35716 1516
rect 35768 1504 35774 1556
rect 36817 1547 36875 1553
rect 36817 1513 36829 1547
rect 36863 1544 36875 1547
rect 37274 1544 37280 1556
rect 36863 1516 37280 1544
rect 36863 1513 36875 1516
rect 36817 1507 36875 1513
rect 37274 1504 37280 1516
rect 37332 1504 37338 1556
rect 37369 1547 37427 1553
rect 37369 1513 37381 1547
rect 37415 1544 37427 1547
rect 39114 1544 39120 1556
rect 37415 1516 39120 1544
rect 37415 1513 37427 1516
rect 37369 1507 37427 1513
rect 39114 1504 39120 1516
rect 39172 1504 39178 1556
rect 39209 1547 39267 1553
rect 39209 1513 39221 1547
rect 39255 1544 39267 1547
rect 41046 1544 41052 1556
rect 39255 1516 41052 1544
rect 39255 1513 39267 1516
rect 39209 1507 39267 1513
rect 41046 1504 41052 1516
rect 41104 1504 41110 1556
rect 41785 1547 41843 1553
rect 41785 1513 41797 1547
rect 41831 1544 41843 1547
rect 43438 1544 43444 1556
rect 41831 1516 43444 1544
rect 41831 1513 41843 1516
rect 41785 1507 41843 1513
rect 43438 1504 43444 1516
rect 43496 1504 43502 1556
rect 43717 1547 43775 1553
rect 43717 1513 43729 1547
rect 43763 1544 43775 1547
rect 44913 1547 44971 1553
rect 43763 1516 44864 1544
rect 43763 1513 43775 1516
rect 43717 1507 43775 1513
rect 33919 1448 35296 1476
rect 35345 1479 35403 1485
rect 33919 1445 33931 1448
rect 33873 1439 33931 1445
rect 35345 1445 35357 1479
rect 35391 1476 35403 1479
rect 37550 1476 37556 1488
rect 35391 1448 37556 1476
rect 35391 1445 35403 1448
rect 35345 1439 35403 1445
rect 37550 1436 37556 1448
rect 37608 1436 37614 1488
rect 37642 1436 37648 1488
rect 37700 1476 37706 1488
rect 37921 1479 37979 1485
rect 37700 1448 37745 1476
rect 37700 1436 37706 1448
rect 37921 1445 37933 1479
rect 37967 1476 37979 1479
rect 39574 1476 39580 1488
rect 37967 1448 39580 1476
rect 37967 1445 37979 1448
rect 37921 1439 37979 1445
rect 39574 1436 39580 1448
rect 39632 1436 39638 1488
rect 40218 1476 40224 1488
rect 40179 1448 40224 1476
rect 40218 1436 40224 1448
rect 40276 1436 40282 1488
rect 40865 1479 40923 1485
rect 40865 1445 40877 1479
rect 40911 1476 40923 1479
rect 42058 1476 42064 1488
rect 40911 1448 42064 1476
rect 40911 1445 40923 1448
rect 40865 1439 40923 1445
rect 42058 1436 42064 1448
rect 42116 1436 42122 1488
rect 42153 1479 42211 1485
rect 42153 1445 42165 1479
rect 42199 1476 42211 1479
rect 42886 1476 42892 1488
rect 42199 1448 42892 1476
rect 42199 1445 42211 1448
rect 42153 1439 42211 1445
rect 42886 1436 42892 1448
rect 42944 1436 42950 1488
rect 42981 1479 43039 1485
rect 42981 1445 42993 1479
rect 43027 1476 43039 1479
rect 44542 1476 44548 1488
rect 43027 1448 44548 1476
rect 43027 1445 43039 1448
rect 42981 1439 43039 1445
rect 44542 1436 44548 1448
rect 44600 1436 44606 1488
rect 44836 1476 44864 1516
rect 44913 1513 44925 1547
rect 44959 1544 44971 1547
rect 46382 1544 46388 1556
rect 44959 1516 46388 1544
rect 44959 1513 44971 1516
rect 44913 1507 44971 1513
rect 46382 1504 46388 1516
rect 46440 1504 46446 1556
rect 46753 1547 46811 1553
rect 46753 1513 46765 1547
rect 46799 1544 46811 1547
rect 48038 1544 48044 1556
rect 46799 1516 48044 1544
rect 46799 1513 46811 1516
rect 46753 1507 46811 1513
rect 48038 1504 48044 1516
rect 48096 1504 48102 1556
rect 48133 1547 48191 1553
rect 48133 1513 48145 1547
rect 48179 1544 48191 1547
rect 49234 1544 49240 1556
rect 48179 1516 49240 1544
rect 48179 1513 48191 1516
rect 48133 1507 48191 1513
rect 49234 1504 49240 1516
rect 49292 1504 49298 1556
rect 49329 1547 49387 1553
rect 49329 1513 49341 1547
rect 49375 1544 49387 1547
rect 49970 1544 49976 1556
rect 49375 1516 49976 1544
rect 49375 1513 49387 1516
rect 49329 1507 49387 1513
rect 49970 1504 49976 1516
rect 50028 1504 50034 1556
rect 50157 1547 50215 1553
rect 50157 1513 50169 1547
rect 50203 1544 50215 1547
rect 51166 1544 51172 1556
rect 50203 1516 51172 1544
rect 50203 1513 50215 1516
rect 50157 1507 50215 1513
rect 51166 1504 51172 1516
rect 51224 1504 51230 1556
rect 51353 1547 51411 1553
rect 51353 1513 51365 1547
rect 51399 1544 51411 1547
rect 52181 1547 52239 1553
rect 51399 1516 52132 1544
rect 51399 1513 51411 1516
rect 51353 1507 51411 1513
rect 45094 1476 45100 1488
rect 44836 1448 45100 1476
rect 45094 1436 45100 1448
rect 45152 1436 45158 1488
rect 45189 1479 45247 1485
rect 45189 1445 45201 1479
rect 45235 1476 45247 1479
rect 46198 1476 46204 1488
rect 45235 1448 46204 1476
rect 45235 1445 45247 1448
rect 45189 1439 45247 1445
rect 46198 1436 46204 1448
rect 46256 1436 46262 1488
rect 47026 1476 47032 1488
rect 46400 1448 47032 1476
rect 33597 1411 33655 1417
rect 33597 1377 33609 1411
rect 33643 1408 33655 1411
rect 35989 1411 36047 1417
rect 33643 1380 35756 1408
rect 33643 1377 33655 1380
rect 33597 1371 33655 1377
rect 34974 1340 34980 1352
rect 33520 1312 34980 1340
rect 34974 1300 34980 1312
rect 35032 1300 35038 1352
rect 35728 1340 35756 1380
rect 35989 1377 36001 1411
rect 36035 1408 36047 1411
rect 37093 1411 37151 1417
rect 36035 1380 37044 1408
rect 36035 1377 36047 1380
rect 35989 1371 36047 1377
rect 36449 1343 36507 1349
rect 35728 1312 35848 1340
rect 35710 1272 35716 1284
rect 33428 1244 35716 1272
rect 35710 1232 35716 1244
rect 35768 1232 35774 1284
rect 34422 1204 34428 1216
rect 31864 1176 34428 1204
rect 34422 1164 34428 1176
rect 34480 1164 34486 1216
rect 35820 1204 35848 1312
rect 36449 1309 36461 1343
rect 36495 1309 36507 1343
rect 37016 1340 37044 1380
rect 37093 1377 37105 1411
rect 37139 1408 37151 1411
rect 38470 1408 38476 1420
rect 37139 1380 38476 1408
rect 37139 1377 37151 1380
rect 37093 1371 37151 1377
rect 38470 1368 38476 1380
rect 38528 1368 38534 1420
rect 38565 1411 38623 1417
rect 38565 1377 38577 1411
rect 38611 1408 38623 1411
rect 39853 1411 39911 1417
rect 38611 1380 39804 1408
rect 38611 1377 38623 1380
rect 38565 1371 38623 1377
rect 38102 1340 38108 1352
rect 37016 1312 38108 1340
rect 36449 1303 36507 1309
rect 36464 1272 36492 1303
rect 38102 1300 38108 1312
rect 38160 1300 38166 1352
rect 38194 1300 38200 1352
rect 38252 1340 38258 1352
rect 38933 1343 38991 1349
rect 38252 1312 38297 1340
rect 38252 1300 38258 1312
rect 38933 1309 38945 1343
rect 38979 1340 38991 1343
rect 39577 1343 39635 1349
rect 38979 1312 39528 1340
rect 38979 1309 38991 1312
rect 38933 1303 38991 1309
rect 38654 1272 38660 1284
rect 36464 1244 38660 1272
rect 38654 1232 38660 1244
rect 38712 1232 38718 1284
rect 36078 1204 36084 1216
rect 35820 1176 36084 1204
rect 36078 1164 36084 1176
rect 36136 1164 36142 1216
rect 39500 1204 39528 1312
rect 39577 1309 39589 1343
rect 39623 1340 39635 1343
rect 39666 1340 39672 1352
rect 39623 1312 39672 1340
rect 39623 1309 39635 1312
rect 39577 1303 39635 1309
rect 39666 1300 39672 1312
rect 39724 1300 39730 1352
rect 39776 1340 39804 1380
rect 39853 1377 39865 1411
rect 39899 1408 39911 1411
rect 40497 1411 40555 1417
rect 39899 1380 40448 1408
rect 39899 1377 39911 1380
rect 39853 1371 39911 1377
rect 40310 1340 40316 1352
rect 39776 1312 40316 1340
rect 40310 1300 40316 1312
rect 40368 1300 40374 1352
rect 40420 1272 40448 1380
rect 40497 1377 40509 1411
rect 40543 1408 40555 1411
rect 41509 1411 41567 1417
rect 40543 1380 41460 1408
rect 40543 1377 40555 1380
rect 40497 1371 40555 1377
rect 41432 1340 41460 1380
rect 41509 1377 41521 1411
rect 41555 1408 41567 1411
rect 42521 1411 42579 1417
rect 41555 1380 42472 1408
rect 41555 1377 41567 1380
rect 41509 1371 41567 1377
rect 42334 1340 42340 1352
rect 41432 1312 42340 1340
rect 42334 1300 42340 1312
rect 42392 1300 42398 1352
rect 42444 1340 42472 1380
rect 42521 1377 42533 1411
rect 42567 1408 42579 1411
rect 44174 1408 44180 1420
rect 42567 1380 44180 1408
rect 42567 1377 42579 1380
rect 42521 1371 42579 1377
rect 44174 1368 44180 1380
rect 44232 1368 44238 1420
rect 44361 1411 44419 1417
rect 44361 1377 44373 1411
rect 44407 1408 44419 1411
rect 44637 1411 44695 1417
rect 44407 1380 44588 1408
rect 44407 1377 44419 1380
rect 44361 1371 44419 1377
rect 43254 1340 43260 1352
rect 42444 1312 43260 1340
rect 43254 1300 43260 1312
rect 43312 1300 43318 1352
rect 43441 1343 43499 1349
rect 43441 1309 43453 1343
rect 43487 1309 43499 1343
rect 43441 1303 43499 1309
rect 41782 1272 41788 1284
rect 40420 1244 41788 1272
rect 41782 1232 41788 1244
rect 41840 1232 41846 1284
rect 40862 1204 40868 1216
rect 39500 1176 40868 1204
rect 40862 1164 40868 1176
rect 40920 1164 40926 1216
rect 43456 1204 43484 1303
rect 44560 1272 44588 1380
rect 44637 1377 44649 1411
rect 44683 1408 44695 1411
rect 45646 1408 45652 1420
rect 44683 1380 45652 1408
rect 44683 1377 44695 1380
rect 44637 1371 44695 1377
rect 45646 1368 45652 1380
rect 45704 1368 45710 1420
rect 45741 1411 45799 1417
rect 45741 1377 45753 1411
rect 45787 1408 45799 1411
rect 46400 1408 46428 1448
rect 47026 1436 47032 1448
rect 47084 1436 47090 1488
rect 47121 1479 47179 1485
rect 47121 1445 47133 1479
rect 47167 1476 47179 1479
rect 48222 1476 48228 1488
rect 47167 1448 48228 1476
rect 47167 1445 47179 1448
rect 47121 1439 47179 1445
rect 48222 1436 48228 1448
rect 48280 1436 48286 1488
rect 48409 1479 48467 1485
rect 48409 1445 48421 1479
rect 48455 1476 48467 1479
rect 48958 1476 48964 1488
rect 48455 1448 48964 1476
rect 48455 1445 48467 1448
rect 48409 1439 48467 1445
rect 48958 1436 48964 1448
rect 49016 1436 49022 1488
rect 50062 1476 50068 1488
rect 49528 1448 50068 1476
rect 45787 1380 46428 1408
rect 46477 1411 46535 1417
rect 45787 1377 45799 1380
rect 45741 1371 45799 1377
rect 46477 1377 46489 1411
rect 46523 1408 46535 1411
rect 47670 1408 47676 1420
rect 46523 1380 47676 1408
rect 46523 1377 46535 1380
rect 46477 1371 46535 1377
rect 47670 1368 47676 1380
rect 47728 1368 47734 1420
rect 47765 1411 47823 1417
rect 47765 1377 47777 1411
rect 47811 1408 47823 1411
rect 48590 1408 48596 1420
rect 47811 1380 48596 1408
rect 47811 1377 47823 1380
rect 47765 1371 47823 1377
rect 48590 1368 48596 1380
rect 48648 1368 48654 1420
rect 48685 1411 48743 1417
rect 48685 1377 48697 1411
rect 48731 1408 48743 1411
rect 49528 1408 49556 1448
rect 50062 1436 50068 1448
rect 50120 1436 50126 1488
rect 50433 1479 50491 1485
rect 50433 1445 50445 1479
rect 50479 1476 50491 1479
rect 51077 1479 51135 1485
rect 50479 1448 50752 1476
rect 50479 1445 50491 1448
rect 50433 1439 50491 1445
rect 48731 1380 48912 1408
rect 48731 1377 48743 1380
rect 48685 1371 48743 1377
rect 45462 1340 45468 1352
rect 45423 1312 45468 1340
rect 45462 1300 45468 1312
rect 45520 1300 45526 1352
rect 46201 1343 46259 1349
rect 46201 1309 46213 1343
rect 46247 1340 46259 1343
rect 47394 1340 47400 1352
rect 46247 1312 47400 1340
rect 46247 1309 46259 1312
rect 46201 1303 46259 1309
rect 47394 1300 47400 1312
rect 47452 1300 47458 1352
rect 47489 1343 47547 1349
rect 47489 1309 47501 1343
rect 47535 1340 47547 1343
rect 48774 1340 48780 1352
rect 47535 1312 48780 1340
rect 47535 1309 47547 1312
rect 47489 1303 47547 1309
rect 48774 1300 48780 1312
rect 48832 1300 48838 1352
rect 45830 1272 45836 1284
rect 44560 1244 45836 1272
rect 45830 1232 45836 1244
rect 45888 1232 45894 1284
rect 48884 1272 48912 1380
rect 48976 1380 49556 1408
rect 49605 1411 49663 1417
rect 48976 1349 49004 1380
rect 49605 1377 49617 1411
rect 49651 1408 49663 1411
rect 50614 1408 50620 1420
rect 49651 1380 50620 1408
rect 49651 1377 49663 1380
rect 49605 1371 49663 1377
rect 50614 1368 50620 1380
rect 50672 1368 50678 1420
rect 48961 1343 49019 1349
rect 48961 1309 48973 1343
rect 49007 1309 49019 1343
rect 50724 1340 50752 1448
rect 51077 1445 51089 1479
rect 51123 1476 51135 1479
rect 51902 1476 51908 1488
rect 51123 1448 51908 1476
rect 51123 1445 51135 1448
rect 51077 1439 51135 1445
rect 51902 1436 51908 1448
rect 51960 1436 51966 1488
rect 52104 1476 52132 1516
rect 52181 1513 52193 1547
rect 52227 1544 52239 1547
rect 53006 1544 53012 1556
rect 52227 1516 53012 1544
rect 52227 1513 52239 1516
rect 52181 1507 52239 1513
rect 53006 1504 53012 1516
rect 53064 1504 53070 1556
rect 55677 1547 55735 1553
rect 55677 1513 55689 1547
rect 55723 1544 55735 1547
rect 55858 1544 55864 1556
rect 55723 1516 55864 1544
rect 55723 1513 55735 1516
rect 55677 1507 55735 1513
rect 55858 1504 55864 1516
rect 55916 1504 55922 1556
rect 55953 1547 56011 1553
rect 55953 1513 55965 1547
rect 55999 1544 56011 1547
rect 56502 1544 56508 1556
rect 55999 1516 56508 1544
rect 55999 1513 56011 1516
rect 55953 1507 56011 1513
rect 56502 1504 56508 1516
rect 56560 1504 56566 1556
rect 56781 1547 56839 1553
rect 56781 1513 56793 1547
rect 56827 1544 56839 1547
rect 58342 1544 58348 1556
rect 56827 1516 58348 1544
rect 56827 1513 56839 1516
rect 56781 1507 56839 1513
rect 58342 1504 58348 1516
rect 58400 1504 58406 1556
rect 52270 1476 52276 1488
rect 52104 1448 52276 1476
rect 52270 1436 52276 1448
rect 52328 1436 52334 1488
rect 52457 1479 52515 1485
rect 52457 1445 52469 1479
rect 52503 1476 52515 1479
rect 52822 1476 52828 1488
rect 52503 1448 52828 1476
rect 52503 1445 52515 1448
rect 52457 1439 52515 1445
rect 52822 1436 52828 1448
rect 52880 1436 52886 1488
rect 53101 1479 53159 1485
rect 53101 1445 53113 1479
rect 53147 1476 53159 1479
rect 53650 1476 53656 1488
rect 53147 1448 53656 1476
rect 53147 1445 53159 1448
rect 53101 1439 53159 1445
rect 53650 1436 53656 1448
rect 53708 1436 53714 1488
rect 53745 1479 53803 1485
rect 53745 1445 53757 1479
rect 53791 1476 53803 1479
rect 54294 1476 54300 1488
rect 53791 1448 54300 1476
rect 53791 1445 53803 1448
rect 53745 1439 53803 1445
rect 54294 1436 54300 1448
rect 54352 1436 54358 1488
rect 54389 1479 54447 1485
rect 54389 1445 54401 1479
rect 54435 1476 54447 1479
rect 54846 1476 54852 1488
rect 54435 1448 54852 1476
rect 54435 1445 54447 1448
rect 54389 1439 54447 1445
rect 54846 1436 54852 1448
rect 54904 1436 54910 1488
rect 55309 1479 55367 1485
rect 55309 1445 55321 1479
rect 55355 1476 55367 1479
rect 56962 1476 56968 1488
rect 55355 1448 56968 1476
rect 55355 1445 55367 1448
rect 55309 1439 55367 1445
rect 56962 1436 56968 1448
rect 57020 1436 57026 1488
rect 57054 1436 57060 1488
rect 57112 1476 57118 1488
rect 57333 1479 57391 1485
rect 57333 1476 57345 1479
rect 57112 1448 57345 1476
rect 57112 1436 57118 1448
rect 57333 1445 57345 1448
rect 57379 1445 57391 1479
rect 57333 1439 57391 1445
rect 57606 1436 57612 1488
rect 57664 1476 57670 1488
rect 57885 1479 57943 1485
rect 57885 1476 57897 1479
rect 57664 1448 57897 1476
rect 57664 1436 57670 1448
rect 57885 1445 57897 1448
rect 57931 1445 57943 1479
rect 57885 1439 57943 1445
rect 50801 1411 50859 1417
rect 50801 1377 50813 1411
rect 50847 1408 50859 1411
rect 51534 1408 51540 1420
rect 50847 1380 51540 1408
rect 50847 1377 50859 1380
rect 50801 1371 50859 1377
rect 51534 1368 51540 1380
rect 51592 1368 51598 1420
rect 51629 1411 51687 1417
rect 51629 1377 51641 1411
rect 51675 1408 51687 1411
rect 53282 1408 53288 1420
rect 51675 1380 52500 1408
rect 51675 1377 51687 1380
rect 51629 1371 51687 1377
rect 52472 1352 52500 1380
rect 52840 1380 53288 1408
rect 51258 1340 51264 1352
rect 50724 1312 51264 1340
rect 48961 1303 49019 1309
rect 51258 1300 51264 1312
rect 51316 1300 51322 1352
rect 52454 1300 52460 1352
rect 52512 1300 52518 1352
rect 52840 1349 52868 1380
rect 53282 1368 53288 1380
rect 53340 1368 53346 1420
rect 53377 1411 53435 1417
rect 53377 1377 53389 1411
rect 53423 1408 53435 1411
rect 53558 1408 53564 1420
rect 53423 1380 53564 1408
rect 53423 1377 53435 1380
rect 53377 1371 53435 1377
rect 53558 1368 53564 1380
rect 53616 1368 53622 1420
rect 54021 1411 54079 1417
rect 54021 1377 54033 1411
rect 54067 1408 54079 1411
rect 54110 1408 54116 1420
rect 54067 1380 54116 1408
rect 54067 1377 54079 1380
rect 54021 1371 54079 1377
rect 54110 1368 54116 1380
rect 54168 1368 54174 1420
rect 54662 1408 54668 1420
rect 54623 1380 54668 1408
rect 54662 1368 54668 1380
rect 54720 1368 54726 1420
rect 54941 1411 54999 1417
rect 54941 1377 54953 1411
rect 54987 1408 54999 1411
rect 55398 1408 55404 1420
rect 54987 1380 55404 1408
rect 54987 1377 54999 1380
rect 54941 1371 54999 1377
rect 55398 1368 55404 1380
rect 55456 1368 55462 1420
rect 56229 1411 56287 1417
rect 56229 1377 56241 1411
rect 56275 1408 56287 1411
rect 56505 1411 56563 1417
rect 56275 1380 56456 1408
rect 56275 1377 56287 1380
rect 56229 1371 56287 1377
rect 52825 1343 52883 1349
rect 52825 1309 52837 1343
rect 52871 1309 52883 1343
rect 56428 1340 56456 1380
rect 56505 1377 56517 1411
rect 56551 1408 56563 1411
rect 56686 1408 56692 1420
rect 56551 1380 56692 1408
rect 56551 1377 56563 1380
rect 56505 1371 56563 1377
rect 56686 1368 56692 1380
rect 56744 1368 56750 1420
rect 57790 1408 57796 1420
rect 57072 1380 57796 1408
rect 56594 1340 56600 1352
rect 56428 1312 56600 1340
rect 52825 1303 52883 1309
rect 56594 1300 56600 1312
rect 56652 1300 56658 1352
rect 57072 1349 57100 1380
rect 57790 1368 57796 1380
rect 57848 1368 57854 1420
rect 57057 1343 57115 1349
rect 57057 1309 57069 1343
rect 57103 1309 57115 1343
rect 57057 1303 57115 1309
rect 57609 1343 57667 1349
rect 57609 1309 57621 1343
rect 57655 1309 57667 1343
rect 57609 1303 57667 1309
rect 49878 1272 49884 1284
rect 48884 1244 49884 1272
rect 49878 1232 49884 1244
rect 49936 1232 49942 1284
rect 56134 1232 56140 1284
rect 56192 1272 56198 1284
rect 57624 1272 57652 1303
rect 56192 1244 57652 1272
rect 56192 1232 56198 1244
rect 45002 1204 45008 1216
rect 43456 1176 45008 1204
rect 45002 1164 45008 1176
rect 45060 1164 45066 1216
rect 1380 1114 58604 1136
rect 1380 1062 3354 1114
rect 3406 1062 19354 1114
rect 19406 1062 35354 1114
rect 35406 1062 51354 1114
rect 51406 1062 58604 1114
rect 1380 1040 58604 1062
<< via1 >>
rect 16764 3612 16816 3664
rect 18880 3612 18932 3664
rect 31576 3544 31628 3596
rect 35164 3544 35216 3596
rect 15108 3476 15160 3528
rect 16764 3476 16816 3528
rect 33232 3476 33284 3528
rect 35900 3476 35952 3528
rect 19340 3408 19392 3460
rect 22560 3408 22612 3460
rect 33784 3408 33836 3460
rect 36084 3408 36136 3460
rect 36176 3408 36228 3460
rect 37004 3408 37056 3460
rect 37280 3408 37332 3460
rect 38292 3408 38344 3460
rect 38844 3408 38896 3460
rect 40684 3408 40736 3460
rect 19892 3340 19944 3392
rect 22192 3340 22244 3392
rect 34520 3340 34572 3392
rect 35532 3340 35584 3392
rect 36912 3340 36964 3392
rect 38752 3340 38804 3392
rect 39120 3340 39172 3392
rect 40868 3340 40920 3392
rect 42800 3340 42852 3392
rect 43260 3340 43312 3392
rect 44272 3340 44324 3392
rect 45100 3340 45152 3392
rect 3354 3238 3406 3290
rect 19354 3238 19406 3290
rect 35354 3238 35406 3290
rect 51354 3238 51406 3290
rect 848 3136 900 3188
rect 5080 3136 5132 3188
rect 13268 3136 13320 3188
rect 14372 3136 14424 3188
rect 1676 3068 1728 3120
rect 3240 3068 3292 3120
rect 7932 3068 7984 3120
rect 2228 3000 2280 3052
rect 2964 3000 3016 3052
rect 3700 3000 3752 3052
rect 4252 3000 4304 3052
rect 4620 3000 4672 3052
rect 5356 3000 5408 3052
rect 5908 3000 5960 3052
rect 6460 3000 6512 3052
rect 7748 3000 7800 3052
rect 9036 3068 9088 3120
rect 8852 3000 8904 3052
rect 12164 3068 12216 3120
rect 10692 3000 10744 3052
rect 11796 3000 11848 3052
rect 13820 3068 13872 3120
rect 15108 3068 15160 3120
rect 14188 3000 14240 3052
rect 17316 3136 17368 3188
rect 19064 3136 19116 3188
rect 19708 3136 19760 3188
rect 16212 3068 16264 3120
rect 16028 3000 16080 3052
rect 18604 3068 18656 3120
rect 18052 3000 18104 3052
rect 20260 3000 20312 3052
rect 21640 3068 21692 3120
rect 22192 3000 22244 3052
rect 22560 3000 22612 3052
rect 24492 3000 24544 3052
rect 25780 3000 25832 3052
rect 27988 3000 28040 3052
rect 28724 3000 28776 3052
rect 31576 3043 31628 3052
rect 31576 3009 31585 3043
rect 31585 3009 31619 3043
rect 31619 3009 31628 3043
rect 31576 3000 31628 3009
rect 34336 3136 34388 3188
rect 32772 3000 32824 3052
rect 34428 3068 34480 3120
rect 33232 3000 33284 3052
rect 33784 3000 33836 3052
rect 36636 3136 36688 3188
rect 38476 3136 38528 3188
rect 38660 3136 38712 3188
rect 39580 3136 39632 3188
rect 37740 3068 37792 3120
rect 37556 3000 37608 3052
rect 2412 2932 2464 2984
rect 3240 2932 3292 2984
rect 4804 2932 4856 2984
rect 6092 2932 6144 2984
rect 6920 2932 6972 2984
rect 7564 2932 7616 2984
rect 9404 2932 9456 2984
rect 10416 2932 10468 2984
rect 11520 2932 11572 2984
rect 2780 2864 2832 2916
rect 1124 2796 1176 2848
rect 3516 2864 3568 2916
rect 7196 2864 7248 2916
rect 8484 2864 8536 2916
rect 9680 2864 9732 2916
rect 11244 2864 11296 2916
rect 5172 2796 5224 2848
rect 5632 2796 5684 2848
rect 7012 2796 7064 2848
rect 9956 2796 10008 2848
rect 11060 2796 11112 2848
rect 12532 2932 12584 2984
rect 13820 2932 13872 2984
rect 14924 2932 14976 2984
rect 16764 2975 16816 2984
rect 16764 2941 16773 2975
rect 16773 2941 16807 2975
rect 16807 2941 16816 2975
rect 16764 2932 16816 2941
rect 18420 2932 18472 2984
rect 20444 2932 20496 2984
rect 22468 2932 22520 2984
rect 13084 2864 13136 2916
rect 15108 2907 15160 2916
rect 15108 2873 15117 2907
rect 15117 2873 15151 2907
rect 15151 2873 15160 2907
rect 15108 2864 15160 2873
rect 15660 2864 15712 2916
rect 17132 2864 17184 2916
rect 18880 2907 18932 2916
rect 18880 2873 18889 2907
rect 18889 2873 18923 2907
rect 18923 2873 18932 2907
rect 18880 2864 18932 2873
rect 18972 2864 19024 2916
rect 20996 2864 21048 2916
rect 12716 2796 12768 2848
rect 14648 2796 14700 2848
rect 16580 2796 16632 2848
rect 19064 2796 19116 2848
rect 19248 2796 19300 2848
rect 20904 2796 20956 2848
rect 29276 2864 29328 2916
rect 32404 2864 32456 2916
rect 35164 2932 35216 2984
rect 37188 2932 37240 2984
rect 25872 2796 25924 2848
rect 34796 2796 34848 2848
rect 35624 2796 35676 2848
rect 35808 2864 35860 2916
rect 36452 2864 36504 2916
rect 36912 2907 36964 2916
rect 36912 2873 36921 2907
rect 36921 2873 36955 2907
rect 36955 2873 36964 2907
rect 39028 3068 39080 3120
rect 39396 3000 39448 3052
rect 39488 3000 39540 3052
rect 42156 3136 42208 3188
rect 42524 3068 42576 3120
rect 40132 2932 40184 2984
rect 41972 3000 42024 3052
rect 42800 3000 42852 3052
rect 44364 3136 44416 3188
rect 44548 3068 44600 3120
rect 44272 3000 44324 3052
rect 46204 3136 46256 3188
rect 46940 3068 46992 3120
rect 46756 3000 46808 3052
rect 48596 3068 48648 3120
rect 48044 3000 48096 3052
rect 48964 3000 49016 3052
rect 50436 3068 50488 3120
rect 50252 3000 50304 3052
rect 51724 3068 51776 3120
rect 51540 3000 51592 3052
rect 52828 3068 52880 3120
rect 53564 3000 53616 3052
rect 54484 3068 54536 3120
rect 54668 3000 54720 3052
rect 55588 3000 55640 3052
rect 58900 3136 58952 3188
rect 41236 2932 41288 2984
rect 43076 2932 43128 2984
rect 45652 2932 45704 2984
rect 47492 2932 47544 2984
rect 49884 2932 49936 2984
rect 50804 2932 50856 2984
rect 52644 2932 52696 2984
rect 53380 2932 53432 2984
rect 55220 2932 55272 2984
rect 58348 3068 58400 3120
rect 56600 3000 56652 3052
rect 58164 3000 58216 3052
rect 56508 2932 56560 2984
rect 36912 2864 36964 2873
rect 36176 2796 36228 2848
rect 37096 2796 37148 2848
rect 39764 2864 39816 2916
rect 41788 2864 41840 2916
rect 43812 2864 43864 2916
rect 44916 2864 44968 2916
rect 47860 2864 47912 2916
rect 49700 2864 49752 2916
rect 50988 2864 51040 2916
rect 52276 2864 52328 2916
rect 53196 2864 53248 2916
rect 54116 2864 54168 2916
rect 55036 2864 55088 2916
rect 56876 2864 56928 2916
rect 57888 2864 57940 2916
rect 38660 2796 38712 2848
rect 38844 2839 38896 2848
rect 38844 2805 38853 2839
rect 38853 2805 38887 2839
rect 38887 2805 38896 2839
rect 38844 2796 38896 2805
rect 39120 2839 39172 2848
rect 39120 2805 39129 2839
rect 39129 2805 39163 2839
rect 39163 2805 39172 2839
rect 39120 2796 39172 2805
rect 39488 2796 39540 2848
rect 41420 2796 41472 2848
rect 44180 2796 44232 2848
rect 45468 2796 45520 2848
rect 47216 2796 47268 2848
rect 49332 2796 49384 2848
rect 59268 2796 59320 2848
rect 11354 2694 11406 2746
rect 27354 2694 27406 2746
rect 43354 2694 43406 2746
rect 1860 2592 1912 2644
rect 3148 2635 3200 2644
rect 3148 2601 3157 2635
rect 3157 2601 3191 2635
rect 3191 2601 3200 2635
rect 3148 2592 3200 2601
rect 4068 2592 4120 2644
rect 8300 2592 8352 2644
rect 10140 2592 10192 2644
rect 11980 2592 12032 2644
rect 15476 2592 15528 2644
rect 17500 2592 17552 2644
rect 21732 2592 21784 2644
rect 22652 2592 22704 2644
rect 23756 2592 23808 2644
rect 23940 2592 23992 2644
rect 24768 2592 24820 2644
rect 25228 2592 25280 2644
rect 25596 2592 25648 2644
rect 25780 2592 25832 2644
rect 26332 2592 26384 2644
rect 26516 2592 26568 2644
rect 27068 2635 27120 2644
rect 27068 2601 27077 2635
rect 27077 2601 27111 2635
rect 27111 2601 27120 2635
rect 27068 2592 27120 2601
rect 27620 2592 27672 2644
rect 28172 2592 28224 2644
rect 29460 2592 29512 2644
rect 30012 2592 30064 2644
rect 30380 2592 30432 2644
rect 30748 2635 30800 2644
rect 30748 2601 30757 2635
rect 30757 2601 30791 2635
rect 30791 2601 30800 2635
rect 30748 2592 30800 2601
rect 31300 2592 31352 2644
rect 33048 2635 33100 2644
rect 33048 2601 33057 2635
rect 33057 2601 33091 2635
rect 33091 2601 33100 2635
rect 33048 2592 33100 2601
rect 33508 2592 33560 2644
rect 34244 2592 34296 2644
rect 37924 2592 37976 2644
rect 40316 2592 40368 2644
rect 43628 2592 43680 2644
rect 46572 2592 46624 2644
rect 48228 2592 48280 2644
rect 50988 2592 51040 2644
rect 52092 2592 52144 2644
rect 53748 2592 53800 2644
rect 55772 2592 55824 2644
rect 56232 2635 56284 2644
rect 56232 2601 56241 2635
rect 56241 2601 56275 2635
rect 56275 2601 56284 2635
rect 56232 2592 56284 2601
rect 57060 2592 57112 2644
rect 572 2524 624 2576
rect 3976 2524 4028 2576
rect 17868 2524 17920 2576
rect 21364 2524 21416 2576
rect 22284 2524 22336 2576
rect 23388 2524 23440 2576
rect 24124 2524 24176 2576
rect 3056 2456 3108 2508
rect 23204 2456 23256 2508
rect 756 2388 808 2440
rect 1308 2320 1360 2372
rect 21548 2388 21600 2440
rect 22928 2388 22980 2440
rect 26056 2524 26108 2576
rect 26148 2524 26200 2576
rect 26424 2524 26476 2576
rect 26884 2524 26936 2576
rect 27528 2524 27580 2576
rect 28908 2524 28960 2576
rect 29828 2524 29880 2576
rect 30564 2524 30616 2576
rect 31668 2524 31720 2576
rect 32956 2524 33008 2576
rect 33692 2524 33744 2576
rect 42708 2524 42760 2576
rect 46020 2524 46072 2576
rect 49148 2524 49200 2576
rect 55956 2524 56008 2576
rect 57612 2524 57664 2576
rect 24676 2456 24728 2508
rect 24768 2456 24820 2508
rect 26240 2456 26292 2508
rect 23112 2320 23164 2372
rect 25504 2388 25556 2440
rect 25596 2388 25648 2440
rect 28264 2456 28316 2508
rect 32220 2456 32272 2508
rect 34060 2456 34112 2508
rect 28356 2388 28408 2440
rect 31852 2388 31904 2440
rect 25044 2320 25096 2372
rect 27804 2320 27856 2372
rect 28448 2320 28500 2372
rect 31300 2320 31352 2372
rect 56048 2388 56100 2440
rect 56324 2456 56376 2508
rect 57428 2388 57480 2440
rect 58716 2320 58768 2372
rect 21088 2252 21140 2304
rect 24952 2252 25004 2304
rect 25320 2252 25372 2304
rect 28540 2252 28592 2304
rect 30380 2252 30432 2304
rect 33140 2252 33192 2304
rect 3354 2150 3406 2202
rect 19354 2150 19406 2202
rect 35354 2150 35406 2202
rect 51354 2150 51406 2202
rect 23848 2048 23900 2100
rect 27068 2048 27120 2100
rect 2044 1912 2096 1964
rect 3700 1955 3752 1964
rect 2596 1844 2648 1896
rect 3700 1921 3709 1955
rect 3709 1921 3743 1955
rect 3743 1921 3752 1955
rect 3700 1912 3752 1921
rect 3976 1955 4028 1964
rect 3976 1921 3985 1955
rect 3985 1921 4019 1955
rect 4019 1921 4028 1955
rect 3976 1912 4028 1921
rect 4160 1912 4212 1964
rect 23296 1980 23348 2032
rect 21088 1955 21140 1964
rect 21088 1921 21097 1955
rect 21097 1921 21131 1955
rect 21131 1921 21140 1955
rect 21088 1912 21140 1921
rect 22008 1912 22060 1964
rect 22836 1912 22888 1964
rect 23112 1955 23164 1964
rect 23112 1921 23121 1955
rect 23121 1921 23155 1955
rect 23155 1921 23164 1955
rect 23112 1912 23164 1921
rect 26148 1980 26200 2032
rect 26332 1980 26384 2032
rect 29460 2048 29512 2100
rect 29552 2048 29604 2100
rect 32404 2048 32456 2100
rect 27712 1980 27764 2032
rect 30656 1980 30708 2032
rect 30932 1980 30984 2032
rect 33692 1980 33744 2032
rect 24768 1912 24820 1964
rect 25044 1955 25096 1964
rect 25044 1921 25053 1955
rect 25053 1921 25087 1955
rect 25087 1921 25096 1955
rect 25044 1912 25096 1921
rect 25320 1955 25372 1964
rect 25320 1921 25329 1955
rect 25329 1921 25363 1955
rect 25363 1921 25372 1955
rect 25320 1912 25372 1921
rect 25596 1955 25648 1964
rect 25596 1921 25605 1955
rect 25605 1921 25639 1955
rect 25639 1921 25648 1955
rect 25596 1912 25648 1921
rect 26608 1912 26660 1964
rect 29644 1912 29696 1964
rect 30380 1955 30432 1964
rect 30380 1921 30389 1955
rect 30389 1921 30423 1955
rect 30423 1921 30432 1955
rect 30380 1912 30432 1921
rect 31116 1955 31168 1964
rect 31116 1921 31125 1955
rect 31125 1921 31159 1955
rect 31159 1921 31168 1955
rect 31116 1912 31168 1921
rect 31392 1912 31444 1964
rect 33324 1912 33376 1964
rect 36268 2048 36320 2100
rect 34152 1980 34204 2032
rect 36636 1980 36688 2032
rect 38200 1980 38252 2032
rect 40132 1980 40184 2032
rect 34796 1912 34848 1964
rect 37188 1912 37240 1964
rect 41420 1912 41472 1964
rect 42064 1912 42116 1964
rect 42708 1912 42760 1964
rect 57980 2048 58032 2100
rect 55864 1980 55916 2032
rect 58532 1980 58584 2032
rect 55680 1955 55732 1964
rect 55680 1921 55689 1955
rect 55689 1921 55723 1955
rect 55723 1921 55732 1955
rect 55680 1912 55732 1921
rect 55956 1955 56008 1964
rect 55956 1921 55965 1955
rect 55965 1921 55999 1955
rect 55999 1921 56008 1955
rect 55956 1912 56008 1921
rect 56232 1955 56284 1964
rect 56232 1921 56241 1955
rect 56241 1921 56275 1955
rect 56275 1921 56284 1955
rect 56232 1912 56284 1921
rect 2780 1776 2832 1828
rect 4252 1844 4304 1896
rect 5080 1887 5132 1896
rect 5080 1853 5089 1887
rect 5089 1853 5123 1887
rect 5123 1853 5132 1887
rect 5080 1844 5132 1853
rect 10324 1844 10376 1896
rect 12716 1844 12768 1896
rect 13268 1844 13320 1896
rect 20628 1844 20680 1896
rect 24400 1844 24452 1896
rect 5172 1776 5224 1828
rect 11060 1776 11112 1828
rect 21180 1776 21232 1828
rect 22008 1776 22060 1828
rect 22836 1776 22888 1828
rect 23572 1776 23624 1828
rect 26240 1776 26292 1828
rect 27252 1776 27304 1828
rect 28816 1776 28868 1828
rect 30840 1844 30892 1896
rect 31576 1844 31628 1896
rect 34244 1844 34296 1896
rect 34428 1844 34480 1896
rect 36820 1844 36872 1896
rect 37280 1844 37332 1896
rect 39028 1844 39080 1896
rect 39672 1844 39724 1896
rect 41604 1844 41656 1896
rect 43996 1844 44048 1896
rect 55220 1844 55272 1896
rect 2872 1751 2924 1760
rect 2872 1717 2881 1751
rect 2881 1717 2915 1751
rect 2915 1717 2924 1751
rect 2872 1708 2924 1717
rect 3240 1708 3292 1760
rect 7196 1708 7248 1760
rect 9588 1708 9640 1760
rect 11612 1708 11664 1760
rect 13452 1708 13504 1760
rect 13820 1751 13872 1760
rect 13820 1717 13829 1751
rect 13829 1717 13863 1751
rect 13863 1717 13872 1751
rect 13820 1708 13872 1717
rect 14556 1708 14608 1760
rect 16948 1708 17000 1760
rect 18236 1708 18288 1760
rect 19524 1708 19576 1760
rect 20352 1708 20404 1760
rect 21732 1708 21784 1760
rect 24308 1708 24360 1760
rect 25964 1708 26016 1760
rect 27896 1708 27948 1760
rect 30748 1776 30800 1828
rect 31484 1776 31536 1828
rect 31760 1776 31812 1828
rect 29092 1708 29144 1760
rect 30012 1708 30064 1760
rect 30564 1708 30616 1760
rect 32036 1708 32088 1760
rect 32220 1776 32272 1828
rect 34704 1776 34756 1828
rect 35072 1776 35124 1828
rect 37372 1776 37424 1828
rect 37648 1776 37700 1828
rect 39764 1776 39816 1828
rect 40224 1776 40276 1828
rect 42156 1776 42208 1828
rect 42892 1776 42944 1828
rect 43812 1776 43864 1828
rect 46572 1776 46624 1828
rect 55956 1776 56008 1828
rect 56784 1819 56836 1828
rect 56784 1785 56793 1819
rect 56793 1785 56827 1819
rect 56827 1785 56836 1819
rect 56784 1776 56836 1785
rect 32772 1708 32824 1760
rect 32864 1708 32916 1760
rect 35164 1708 35216 1760
rect 35716 1708 35768 1760
rect 37832 1708 37884 1760
rect 39948 1708 40000 1760
rect 42800 1708 42852 1760
rect 44732 1708 44784 1760
rect 45468 1708 45520 1760
rect 46940 1708 46992 1760
rect 49516 1708 49568 1760
rect 50988 1708 51040 1760
rect 55588 1708 55640 1760
rect 56508 1751 56560 1760
rect 56508 1717 56517 1751
rect 56517 1717 56551 1751
rect 56551 1717 56560 1751
rect 56508 1708 56560 1717
rect 56600 1708 56652 1760
rect 58900 1776 58952 1828
rect 59084 1708 59136 1760
rect 11354 1606 11406 1658
rect 27354 1606 27406 1658
rect 43354 1606 43406 1658
rect 572 1504 624 1556
rect 3884 1504 3936 1556
rect 6644 1504 6696 1556
rect 8116 1504 8168 1556
rect 1492 1436 1544 1488
rect 1308 1368 1360 1420
rect 1860 1368 1912 1420
rect 2412 1368 2464 1420
rect 3700 1436 3752 1488
rect 4804 1436 4856 1488
rect 5724 1436 5776 1488
rect 6368 1436 6420 1488
rect 7380 1436 7432 1488
rect 8484 1504 8536 1556
rect 9772 1504 9824 1556
rect 11520 1504 11572 1556
rect 14004 1504 14056 1556
rect 18788 1504 18840 1556
rect 20076 1504 20128 1556
rect 22928 1547 22980 1556
rect 22928 1513 22937 1547
rect 22937 1513 22971 1547
rect 22971 1513 22980 1547
rect 22928 1504 22980 1513
rect 23020 1504 23072 1556
rect 25044 1504 25096 1556
rect 27620 1504 27672 1556
rect 27712 1547 27764 1556
rect 27712 1513 27721 1547
rect 27721 1513 27755 1547
rect 27755 1513 27764 1547
rect 27712 1504 27764 1513
rect 28448 1504 28500 1556
rect 9220 1436 9272 1488
rect 10876 1436 10928 1488
rect 12164 1436 12216 1488
rect 16212 1436 16264 1488
rect 17684 1436 17736 1488
rect 18604 1436 18656 1488
rect 19892 1436 19944 1488
rect 3240 1368 3292 1420
rect 3516 1368 3568 1420
rect 940 1232 992 1284
rect 4436 1368 4488 1420
rect 4988 1368 5040 1420
rect 5540 1368 5592 1420
rect 6092 1368 6144 1420
rect 6828 1368 6880 1420
rect 7932 1368 7984 1420
rect 8852 1368 8904 1420
rect 9956 1368 10008 1420
rect 7656 1300 7708 1352
rect 9036 1300 9088 1352
rect 10600 1300 10652 1352
rect 11980 1368 12032 1420
rect 12348 1368 12400 1420
rect 12900 1411 12952 1420
rect 12900 1377 12909 1411
rect 12909 1377 12943 1411
rect 12943 1377 12952 1411
rect 12900 1368 12952 1377
rect 14188 1368 14240 1420
rect 14740 1368 14792 1420
rect 15108 1368 15160 1420
rect 15292 1411 15344 1420
rect 15292 1377 15301 1411
rect 15301 1377 15335 1411
rect 15335 1377 15344 1411
rect 15292 1368 15344 1377
rect 15660 1368 15712 1420
rect 15844 1368 15896 1420
rect 16396 1411 16448 1420
rect 16396 1377 16405 1411
rect 16405 1377 16439 1411
rect 16439 1377 16448 1411
rect 16396 1368 16448 1377
rect 16580 1368 16632 1420
rect 17132 1368 17184 1420
rect 17500 1368 17552 1420
rect 18144 1368 18196 1420
rect 18972 1368 19024 1420
rect 19524 1368 19576 1420
rect 20352 1411 20404 1420
rect 20352 1377 20361 1411
rect 20361 1377 20395 1411
rect 20395 1377 20404 1411
rect 20352 1368 20404 1377
rect 20444 1368 20496 1420
rect 22284 1436 22336 1488
rect 23756 1436 23808 1488
rect 20996 1368 21048 1420
rect 24768 1436 24820 1488
rect 26332 1479 26384 1488
rect 26332 1445 26341 1479
rect 26341 1445 26375 1479
rect 26375 1445 26384 1479
rect 26332 1436 26384 1445
rect 26608 1479 26660 1488
rect 26608 1445 26617 1479
rect 26617 1445 26651 1479
rect 26651 1445 26660 1479
rect 26608 1436 26660 1445
rect 29092 1504 29144 1556
rect 30564 1504 30616 1556
rect 31392 1504 31444 1556
rect 31576 1547 31628 1556
rect 31576 1513 31585 1547
rect 31585 1513 31619 1547
rect 31619 1513 31628 1547
rect 31576 1504 31628 1513
rect 32220 1547 32272 1556
rect 32220 1513 32229 1547
rect 32229 1513 32263 1547
rect 32263 1513 32272 1547
rect 32220 1504 32272 1513
rect 30748 1436 30800 1488
rect 30932 1479 30984 1488
rect 30932 1445 30941 1479
rect 30941 1445 30975 1479
rect 30975 1445 30984 1479
rect 30932 1436 30984 1445
rect 33784 1504 33836 1556
rect 34152 1547 34204 1556
rect 34152 1513 34161 1547
rect 34161 1513 34195 1547
rect 34195 1513 34204 1547
rect 34152 1504 34204 1513
rect 34428 1547 34480 1556
rect 34428 1513 34437 1547
rect 34437 1513 34471 1547
rect 34471 1513 34480 1547
rect 34428 1504 34480 1513
rect 34796 1547 34848 1556
rect 34796 1513 34805 1547
rect 34805 1513 34839 1547
rect 34839 1513 34848 1547
rect 34796 1504 34848 1513
rect 35072 1547 35124 1556
rect 35072 1513 35081 1547
rect 35081 1513 35115 1547
rect 35115 1513 35124 1547
rect 35072 1504 35124 1513
rect 23388 1300 23440 1352
rect 23848 1300 23900 1352
rect 25780 1232 25832 1284
rect 25412 1164 25464 1216
rect 26148 1164 26200 1216
rect 26700 1164 26752 1216
rect 30196 1368 30248 1420
rect 32588 1368 32640 1420
rect 32864 1411 32916 1420
rect 32864 1377 32873 1411
rect 32873 1377 32907 1411
rect 32907 1377 32916 1411
rect 32864 1368 32916 1377
rect 29552 1343 29604 1352
rect 28816 1232 28868 1284
rect 29552 1309 29561 1343
rect 29561 1309 29595 1343
rect 29595 1309 29604 1343
rect 29552 1300 29604 1309
rect 31760 1300 31812 1352
rect 30380 1164 30432 1216
rect 31760 1164 31812 1216
rect 35532 1504 35584 1556
rect 35716 1547 35768 1556
rect 35716 1513 35725 1547
rect 35725 1513 35759 1547
rect 35759 1513 35768 1547
rect 35716 1504 35768 1513
rect 37280 1504 37332 1556
rect 39120 1504 39172 1556
rect 41052 1504 41104 1556
rect 43444 1504 43496 1556
rect 37556 1436 37608 1488
rect 37648 1479 37700 1488
rect 37648 1445 37657 1479
rect 37657 1445 37691 1479
rect 37691 1445 37700 1479
rect 37648 1436 37700 1445
rect 39580 1436 39632 1488
rect 40224 1479 40276 1488
rect 40224 1445 40233 1479
rect 40233 1445 40267 1479
rect 40267 1445 40276 1479
rect 40224 1436 40276 1445
rect 42064 1436 42116 1488
rect 42892 1436 42944 1488
rect 44548 1436 44600 1488
rect 46388 1504 46440 1556
rect 48044 1504 48096 1556
rect 49240 1504 49292 1556
rect 49976 1504 50028 1556
rect 51172 1504 51224 1556
rect 45100 1436 45152 1488
rect 46204 1436 46256 1488
rect 34980 1300 35032 1352
rect 35716 1232 35768 1284
rect 34428 1164 34480 1216
rect 38476 1368 38528 1420
rect 38108 1300 38160 1352
rect 38200 1343 38252 1352
rect 38200 1309 38209 1343
rect 38209 1309 38243 1343
rect 38243 1309 38252 1343
rect 38200 1300 38252 1309
rect 38660 1232 38712 1284
rect 36084 1164 36136 1216
rect 39672 1300 39724 1352
rect 40316 1300 40368 1352
rect 42340 1300 42392 1352
rect 44180 1368 44232 1420
rect 43260 1300 43312 1352
rect 41788 1232 41840 1284
rect 40868 1164 40920 1216
rect 45652 1368 45704 1420
rect 47032 1436 47084 1488
rect 48228 1436 48280 1488
rect 48964 1436 49016 1488
rect 47676 1368 47728 1420
rect 48596 1368 48648 1420
rect 50068 1436 50120 1488
rect 45468 1343 45520 1352
rect 45468 1309 45477 1343
rect 45477 1309 45511 1343
rect 45511 1309 45520 1343
rect 45468 1300 45520 1309
rect 47400 1300 47452 1352
rect 48780 1300 48832 1352
rect 45836 1232 45888 1284
rect 50620 1368 50672 1420
rect 51908 1436 51960 1488
rect 53012 1504 53064 1556
rect 55864 1504 55916 1556
rect 56508 1504 56560 1556
rect 58348 1504 58400 1556
rect 52276 1436 52328 1488
rect 52828 1436 52880 1488
rect 53656 1436 53708 1488
rect 54300 1436 54352 1488
rect 54852 1436 54904 1488
rect 56968 1436 57020 1488
rect 57060 1436 57112 1488
rect 57612 1436 57664 1488
rect 51540 1368 51592 1420
rect 51264 1300 51316 1352
rect 52460 1300 52512 1352
rect 53288 1368 53340 1420
rect 53564 1368 53616 1420
rect 54116 1368 54168 1420
rect 54668 1411 54720 1420
rect 54668 1377 54677 1411
rect 54677 1377 54711 1411
rect 54711 1377 54720 1411
rect 54668 1368 54720 1377
rect 55404 1368 55456 1420
rect 56692 1368 56744 1420
rect 56600 1300 56652 1352
rect 57796 1368 57848 1420
rect 49884 1232 49936 1284
rect 56140 1232 56192 1284
rect 45008 1164 45060 1216
rect 3354 1062 3406 1114
rect 19354 1062 19406 1114
rect 35354 1062 35406 1114
rect 51354 1062 51406 1114
<< metal2 >>
rect 570 3800 626 4600
rect 754 3800 810 4600
rect 1122 3800 1178 4600
rect 1306 3800 1362 4600
rect 1674 3800 1730 4600
rect 1858 3800 1914 4600
rect 2226 3800 2282 4600
rect 2410 3800 2466 4600
rect 2778 3800 2834 4600
rect 2962 3800 3018 4600
rect 3146 3800 3202 4600
rect 3514 3800 3570 4600
rect 3698 3800 3754 4600
rect 4066 3800 4122 4600
rect 4250 3800 4306 4600
rect 4618 3800 4674 4600
rect 4802 3800 4858 4600
rect 5170 3800 5226 4600
rect 5354 3800 5410 4600
rect 5538 3800 5594 4600
rect 5906 3800 5962 4600
rect 6090 3800 6146 4600
rect 6458 3800 6514 4600
rect 6642 3800 6698 4600
rect 7010 3800 7066 4600
rect 7194 3800 7250 4600
rect 7562 3800 7618 4600
rect 7746 3800 7802 4600
rect 7930 3800 7986 4600
rect 8298 3800 8354 4600
rect 8482 3800 8538 4600
rect 8850 3800 8906 4600
rect 9034 3800 9090 4600
rect 9402 3800 9458 4600
rect 9586 3800 9642 4600
rect 9954 3800 10010 4600
rect 10138 3800 10194 4600
rect 10322 3800 10378 4600
rect 10690 3800 10746 4600
rect 10874 3800 10930 4600
rect 11242 3800 11298 4600
rect 11426 3800 11482 4600
rect 11794 3800 11850 4600
rect 11978 3800 12034 4600
rect 12162 3800 12218 4600
rect 12530 3800 12586 4600
rect 12714 3800 12770 4600
rect 13082 3800 13138 4600
rect 13266 3800 13322 4600
rect 13634 3800 13690 4600
rect 13818 3800 13874 4600
rect 14186 3800 14242 4600
rect 14370 3800 14426 4600
rect 14554 3800 14610 4600
rect 14922 3800 14978 4600
rect 15106 3800 15162 4600
rect 15474 3800 15530 4600
rect 15658 3800 15714 4600
rect 16026 3800 16082 4600
rect 16210 3800 16266 4600
rect 16578 3800 16634 4600
rect 16762 3800 16818 4600
rect 16946 3800 17002 4600
rect 17314 3800 17370 4600
rect 17498 3800 17554 4600
rect 17866 3800 17922 4600
rect 18050 3800 18106 4600
rect 18418 3800 18474 4600
rect 18602 3800 18658 4600
rect 18970 3800 19026 4600
rect 19154 3800 19210 4600
rect 19338 3800 19394 4600
rect 19706 3800 19762 4600
rect 19890 3800 19946 4600
rect 20258 3800 20314 4600
rect 20442 3800 20498 4600
rect 20810 3800 20866 4600
rect 20994 3800 21050 4600
rect 21362 3800 21418 4600
rect 21546 3800 21602 4600
rect 21730 3800 21786 4600
rect 22098 3800 22154 4600
rect 22282 3800 22338 4600
rect 22650 3800 22706 4600
rect 22834 3800 22890 4600
rect 23202 3800 23258 4600
rect 23386 3800 23442 4600
rect 23754 3800 23810 4600
rect 23938 3800 23994 4600
rect 24122 3800 24178 4600
rect 24490 3800 24546 4600
rect 24674 3800 24730 4600
rect 25042 3800 25098 4600
rect 25226 3800 25282 4600
rect 25594 3800 25650 4600
rect 25778 3800 25834 4600
rect 25962 3800 26018 4600
rect 26330 3800 26386 4600
rect 26514 3800 26570 4600
rect 26882 3800 26938 4600
rect 27066 3800 27122 4600
rect 27434 3800 27490 4600
rect 27618 3800 27674 4600
rect 27986 3800 28042 4600
rect 28170 3800 28226 4600
rect 28354 3800 28410 4600
rect 28722 3800 28778 4600
rect 28906 3800 28962 4600
rect 29274 3800 29330 4600
rect 29458 3800 29514 4600
rect 29826 3800 29882 4600
rect 30010 3800 30066 4600
rect 30378 3800 30434 4600
rect 30562 3800 30618 4600
rect 30746 3800 30802 4600
rect 31114 3800 31170 4600
rect 31298 3800 31354 4600
rect 31666 3800 31722 4600
rect 31850 3800 31906 4600
rect 32218 3800 32274 4600
rect 32402 3800 32458 4600
rect 32770 3800 32826 4600
rect 32954 3800 33010 4600
rect 33138 3800 33194 4600
rect 33506 3800 33562 4600
rect 33690 3800 33746 4600
rect 34058 3800 34114 4600
rect 34242 3800 34298 4600
rect 34610 3800 34666 4600
rect 34794 3800 34850 4600
rect 35162 3800 35218 4600
rect 35346 3800 35402 4600
rect 35530 3800 35586 4600
rect 35898 3800 35954 4600
rect 36082 3800 36138 4600
rect 36450 3800 36506 4600
rect 36634 3800 36690 4600
rect 37002 3800 37058 4600
rect 37186 3800 37242 4600
rect 37554 3800 37610 4600
rect 37738 3800 37794 4600
rect 37922 3800 37978 4600
rect 38290 3800 38346 4600
rect 38474 3800 38530 4600
rect 38842 3800 38898 4600
rect 39026 3800 39082 4600
rect 39394 3800 39450 4600
rect 39578 3800 39634 4600
rect 39762 3800 39818 4600
rect 40130 3800 40186 4600
rect 40314 3800 40370 4600
rect 40682 3800 40738 4600
rect 40866 3800 40922 4600
rect 41234 3800 41290 4600
rect 41418 3800 41474 4600
rect 41786 3800 41842 4600
rect 41970 3800 42026 4600
rect 42154 3800 42210 4600
rect 42522 3800 42578 4600
rect 42706 3800 42762 4600
rect 43074 3800 43130 4600
rect 43258 3800 43314 4600
rect 43626 3800 43682 4600
rect 43810 3800 43866 4600
rect 44178 3800 44234 4600
rect 44362 3800 44418 4600
rect 44546 3800 44602 4600
rect 44914 3800 44970 4600
rect 45098 3800 45154 4600
rect 45466 3800 45522 4600
rect 45650 3800 45706 4600
rect 46018 3800 46074 4600
rect 46202 3800 46258 4600
rect 46570 3800 46626 4600
rect 46754 3800 46810 4600
rect 46938 3800 46994 4600
rect 47306 3800 47362 4600
rect 47490 3800 47546 4600
rect 47858 3800 47914 4600
rect 48042 3800 48098 4600
rect 48410 3800 48466 4600
rect 48594 3800 48650 4600
rect 48962 3800 49018 4600
rect 49146 3800 49202 4600
rect 49330 3800 49386 4600
rect 49698 3800 49754 4600
rect 49882 3800 49938 4600
rect 50250 3800 50306 4600
rect 50434 3800 50490 4600
rect 50802 3800 50858 4600
rect 50986 3800 51042 4600
rect 51354 3800 51410 4600
rect 51538 3800 51594 4600
rect 51722 3800 51778 4600
rect 52090 3800 52146 4600
rect 52274 3800 52330 4600
rect 52642 3800 52698 4600
rect 52826 3800 52882 4600
rect 53194 3800 53250 4600
rect 53378 3800 53434 4600
rect 53562 3800 53618 4600
rect 53930 3800 53986 4600
rect 54114 3800 54170 4600
rect 54482 3800 54538 4600
rect 54666 3800 54722 4600
rect 55034 3800 55090 4600
rect 55218 3800 55274 4600
rect 55586 3800 55642 4600
rect 55770 3800 55826 4600
rect 55954 3800 56010 4600
rect 56322 3800 56378 4600
rect 56506 3800 56562 4600
rect 56874 3800 56930 4600
rect 57058 3800 57114 4600
rect 57426 3800 57482 4600
rect 57610 3800 57666 4600
rect 57978 3800 58034 4600
rect 58162 3800 58218 4600
rect 58346 3800 58402 4600
rect 58714 3800 58770 4600
rect 58898 3800 58954 4600
rect 59266 3800 59322 4600
rect 584 2582 612 3800
rect 572 2576 624 2582
rect 572 2518 624 2524
rect 768 2446 796 3800
rect 848 3188 900 3194
rect 848 3130 900 3136
rect 756 2440 808 2446
rect 756 2382 808 2388
rect 572 1556 624 1562
rect 572 1498 624 1504
rect 584 800 612 1498
rect 860 898 888 3130
rect 1136 2854 1164 3800
rect 1124 2848 1176 2854
rect 1124 2790 1176 2796
rect 1320 2378 1348 3800
rect 1688 3126 1716 3800
rect 1676 3120 1728 3126
rect 1676 3062 1728 3068
rect 1872 2650 1900 3800
rect 2240 3058 2268 3800
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 2424 2990 2452 3800
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 2792 2922 2820 3800
rect 2976 3058 3004 3800
rect 3160 3754 3188 3800
rect 3068 3726 3188 3754
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 2780 2916 2832 2922
rect 2780 2858 2832 2864
rect 1860 2644 1912 2650
rect 1860 2586 1912 2592
rect 3068 2514 3096 3726
rect 3146 3632 3202 3641
rect 3146 3567 3202 3576
rect 3160 2650 3188 3567
rect 3350 3290 3410 3312
rect 3350 3238 3354 3290
rect 3406 3238 3410 3290
rect 3240 3120 3292 3126
rect 3240 3062 3292 3068
rect 3252 2990 3280 3062
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 1308 2372 1360 2378
rect 1308 2314 1360 2320
rect 3350 2202 3410 3238
rect 3528 2922 3556 3800
rect 3712 3058 3740 3800
rect 3974 3088 4030 3097
rect 3700 3052 3752 3058
rect 3974 3023 4030 3032
rect 3700 2994 3752 3000
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 3988 2582 4016 3023
rect 4080 2650 4108 3800
rect 4264 3058 4292 3800
rect 4632 3058 4660 3800
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4816 2990 4844 3800
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 4158 2816 4214 2825
rect 4158 2751 4214 2760
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 3976 2576 4028 2582
rect 3976 2518 4028 2524
rect 3350 2150 3354 2202
rect 3406 2150 3410 2202
rect 2044 1964 2096 1970
rect 2044 1906 2096 1912
rect 1492 1488 1544 1494
rect 1492 1430 1544 1436
rect 1308 1420 1360 1426
rect 1308 1362 1360 1368
rect 940 1284 992 1290
rect 940 1226 992 1232
rect 768 870 888 898
rect 768 800 796 870
rect 952 800 980 1226
rect 1320 800 1348 1362
rect 1504 800 1532 1430
rect 1860 1420 1912 1426
rect 1860 1362 1912 1368
rect 1872 800 1900 1362
rect 2056 800 2084 1906
rect 2596 1896 2648 1902
rect 2596 1838 2648 1844
rect 2412 1420 2464 1426
rect 2412 1362 2464 1368
rect 2424 800 2452 1362
rect 2608 800 2636 1838
rect 2780 1828 2832 1834
rect 2780 1770 2832 1776
rect 2792 800 2820 1770
rect 2872 1760 2924 1766
rect 3240 1760 3292 1766
rect 2872 1702 2924 1708
rect 3160 1720 3240 1748
rect 2884 1057 2912 1702
rect 2870 1048 2926 1057
rect 2870 983 2926 992
rect 3160 800 3188 1720
rect 3240 1702 3292 1708
rect 3240 1420 3292 1426
rect 3240 1362 3292 1368
rect 3252 898 3280 1362
rect 3350 1268 3410 2150
rect 3974 2136 4030 2145
rect 3974 2071 4030 2080
rect 3698 2000 3754 2009
rect 3988 1970 4016 2071
rect 4172 1970 4200 2751
rect 3698 1935 3700 1944
rect 3752 1935 3754 1944
rect 3976 1964 4028 1970
rect 3700 1906 3752 1912
rect 3976 1906 4028 1912
rect 4160 1964 4212 1970
rect 4160 1906 4212 1912
rect 5092 1902 5120 3130
rect 5184 2854 5212 3800
rect 5368 3058 5396 3800
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5172 2848 5224 2854
rect 5552 2836 5580 3800
rect 5920 3058 5948 3800
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 6104 2990 6132 3800
rect 6472 3058 6500 3800
rect 6656 3074 6684 3800
rect 6460 3052 6512 3058
rect 6656 3046 6960 3074
rect 6460 2994 6512 3000
rect 6932 2990 6960 3046
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 7024 2854 7052 3800
rect 7208 2922 7236 3800
rect 7576 2990 7604 3800
rect 7760 3058 7788 3800
rect 7944 3126 7972 3800
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7564 2984 7616 2990
rect 7564 2926 7616 2932
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 5632 2848 5684 2854
rect 5552 2808 5632 2836
rect 5172 2790 5224 2796
rect 5632 2790 5684 2796
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 8312 2650 8340 3800
rect 8496 2922 8524 3800
rect 8864 3058 8892 3800
rect 9048 3126 9076 3800
rect 9036 3120 9088 3126
rect 9036 3062 9088 3068
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 9416 2990 9444 3800
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9600 2938 9628 3800
rect 9600 2922 9720 2938
rect 8484 2916 8536 2922
rect 9600 2916 9732 2922
rect 9600 2910 9680 2916
rect 8484 2858 8536 2864
rect 9680 2858 9732 2864
rect 9968 2854 9996 3800
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 10152 2650 10180 3800
rect 10336 2972 10364 3800
rect 10704 3058 10732 3800
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10416 2984 10468 2990
rect 10336 2944 10416 2972
rect 10416 2926 10468 2932
rect 10888 2836 10916 3800
rect 11256 2922 11284 3800
rect 11244 2916 11296 2922
rect 11244 2858 11296 2864
rect 11060 2848 11112 2854
rect 10888 2808 11060 2836
rect 11060 2790 11112 2796
rect 11350 2746 11410 3312
rect 11440 2972 11468 3800
rect 11808 3058 11836 3800
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11520 2984 11572 2990
rect 11440 2944 11520 2972
rect 11520 2926 11572 2932
rect 11350 2694 11354 2746
rect 11406 2694 11410 2746
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 11350 2348 11410 2694
rect 11992 2650 12020 3800
rect 12176 3126 12204 3800
rect 12164 3120 12216 3126
rect 12164 3062 12216 3068
rect 12544 2990 12572 3800
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 12728 2854 12756 3800
rect 13096 2922 13124 3800
rect 13280 3194 13308 3800
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13648 2972 13676 3800
rect 13832 3126 13860 3800
rect 13820 3120 13872 3126
rect 13820 3062 13872 3068
rect 14200 3058 14228 3800
rect 14384 3194 14412 3800
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 13820 2984 13872 2990
rect 13648 2944 13820 2972
rect 13820 2926 13872 2932
rect 13084 2916 13136 2922
rect 13084 2858 13136 2864
rect 12716 2848 12768 2854
rect 14568 2836 14596 3800
rect 14936 2990 14964 3800
rect 15120 3534 15148 3800
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 15108 3120 15160 3126
rect 15108 3062 15160 3068
rect 14924 2984 14976 2990
rect 14924 2926 14976 2932
rect 15120 2922 15148 3062
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 14648 2848 14700 2854
rect 14568 2808 14648 2836
rect 12716 2790 12768 2796
rect 14648 2790 14700 2796
rect 15488 2650 15516 3800
rect 15672 2922 15700 3800
rect 16040 3058 16068 3800
rect 16224 3126 16252 3800
rect 16212 3120 16264 3126
rect 16212 3062 16264 3068
rect 16028 3052 16080 3058
rect 16028 2994 16080 3000
rect 15660 2916 15712 2922
rect 15660 2858 15712 2864
rect 16592 2854 16620 3800
rect 16776 3670 16804 3800
rect 16764 3664 16816 3670
rect 16764 3606 16816 3612
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16776 2990 16804 3470
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16960 2938 16988 3800
rect 17328 3194 17356 3800
rect 17316 3188 17368 3194
rect 17316 3130 17368 3136
rect 16960 2922 17172 2938
rect 16960 2916 17184 2922
rect 16960 2910 17132 2916
rect 17132 2858 17184 2864
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 17512 2650 17540 3800
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 17880 2582 17908 3800
rect 18064 3058 18092 3800
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 18432 2990 18460 3800
rect 18616 3126 18644 3800
rect 18880 3664 18932 3670
rect 18880 3606 18932 3612
rect 18604 3120 18656 3126
rect 18604 3062 18656 3068
rect 18420 2984 18472 2990
rect 18420 2926 18472 2932
rect 18892 2922 18920 3606
rect 18984 2922 19012 3800
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 18880 2916 18932 2922
rect 18880 2858 18932 2864
rect 18972 2916 19024 2922
rect 18972 2858 19024 2864
rect 19076 2854 19104 3130
rect 19168 2938 19196 3800
rect 19352 3466 19380 3800
rect 19340 3460 19392 3466
rect 19340 3402 19392 3408
rect 19350 3290 19410 3312
rect 19350 3238 19354 3290
rect 19406 3238 19410 3290
rect 19168 2910 19288 2938
rect 19260 2854 19288 2910
rect 19064 2848 19116 2854
rect 19064 2790 19116 2796
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 17868 2576 17920 2582
rect 17868 2518 17920 2524
rect 11350 2292 11352 2348
rect 11408 2292 11410 2348
rect 4252 1896 4304 1902
rect 4252 1838 4304 1844
rect 5080 1896 5132 1902
rect 5080 1838 5132 1844
rect 10324 1896 10376 1902
rect 10324 1838 10376 1844
rect 3884 1556 3936 1562
rect 3884 1498 3936 1504
rect 3700 1488 3752 1494
rect 3514 1456 3570 1465
rect 3700 1430 3752 1436
rect 3514 1391 3516 1400
rect 3568 1391 3570 1400
rect 3516 1362 3568 1368
rect 3350 1212 3352 1268
rect 3408 1212 3410 1268
rect 3350 1114 3410 1212
rect 3350 1062 3354 1114
rect 3406 1062 3410 1114
rect 3350 1040 3410 1062
rect 3252 870 3372 898
rect 3344 800 3372 870
rect 3712 800 3740 1430
rect 3896 800 3924 1498
rect 4264 800 4292 1838
rect 5172 1828 5224 1834
rect 5172 1770 5224 1776
rect 4804 1488 4856 1494
rect 4804 1430 4856 1436
rect 4436 1420 4488 1426
rect 4436 1362 4488 1368
rect 4448 800 4476 1362
rect 4816 800 4844 1430
rect 4988 1420 5040 1426
rect 4988 1362 5040 1368
rect 5000 800 5028 1362
rect 5184 800 5212 1770
rect 7196 1760 7248 1766
rect 7196 1702 7248 1708
rect 9588 1760 9640 1766
rect 9588 1702 9640 1708
rect 6644 1556 6696 1562
rect 6644 1498 6696 1504
rect 5724 1488 5776 1494
rect 5724 1430 5776 1436
rect 6368 1488 6420 1494
rect 6368 1430 6420 1436
rect 5540 1420 5592 1426
rect 5540 1362 5592 1368
rect 5552 800 5580 1362
rect 5736 800 5764 1430
rect 6092 1420 6144 1426
rect 6092 1362 6144 1368
rect 6104 800 6132 1362
rect 6380 898 6408 1430
rect 6288 870 6408 898
rect 6288 800 6316 870
rect 6656 800 6684 1498
rect 6828 1420 6880 1426
rect 6828 1362 6880 1368
rect 6840 800 6868 1362
rect 7208 800 7236 1702
rect 8116 1556 8168 1562
rect 8116 1498 8168 1504
rect 8484 1556 8536 1562
rect 8484 1498 8536 1504
rect 7380 1488 7432 1494
rect 7380 1430 7432 1436
rect 7392 800 7420 1430
rect 7932 1420 7984 1426
rect 7932 1362 7984 1368
rect 7656 1352 7708 1358
rect 7656 1294 7708 1300
rect 7668 898 7696 1294
rect 7576 870 7696 898
rect 7576 800 7604 870
rect 7944 800 7972 1362
rect 8128 800 8156 1498
rect 8496 800 8524 1498
rect 9220 1488 9272 1494
rect 9220 1430 9272 1436
rect 8852 1420 8904 1426
rect 8680 1380 8852 1408
rect 8680 800 8708 1380
rect 8852 1362 8904 1368
rect 9036 1352 9088 1358
rect 9036 1294 9088 1300
rect 9048 800 9076 1294
rect 9232 800 9260 1430
rect 9600 800 9628 1702
rect 9772 1556 9824 1562
rect 9772 1498 9824 1504
rect 9784 800 9812 1498
rect 9956 1420 10008 1426
rect 9956 1362 10008 1368
rect 9968 800 9996 1362
rect 10336 800 10364 1838
rect 11060 1828 11112 1834
rect 11060 1770 11112 1776
rect 10876 1488 10928 1494
rect 10876 1430 10928 1436
rect 10600 1352 10652 1358
rect 10600 1294 10652 1300
rect 10612 898 10640 1294
rect 10520 870 10640 898
rect 10520 800 10548 870
rect 10888 800 10916 1430
rect 11072 800 11100 1770
rect 11350 1658 11410 2292
rect 19350 2202 19410 3238
rect 19720 3194 19748 3800
rect 19904 3398 19932 3800
rect 19892 3392 19944 3398
rect 19892 3334 19944 3340
rect 19708 3188 19760 3194
rect 19708 3130 19760 3136
rect 20272 3058 20300 3800
rect 20260 3052 20312 3058
rect 20260 2994 20312 3000
rect 20456 2990 20484 3800
rect 20444 2984 20496 2990
rect 20444 2926 20496 2932
rect 20824 2938 20852 3800
rect 20824 2910 20944 2938
rect 21008 2922 21036 3800
rect 20916 2854 20944 2910
rect 20996 2916 21048 2922
rect 20996 2858 21048 2864
rect 20904 2848 20956 2854
rect 20904 2790 20956 2796
rect 21376 2582 21404 3800
rect 21364 2576 21416 2582
rect 21364 2518 21416 2524
rect 21560 2446 21588 3800
rect 21640 3120 21692 3126
rect 21640 3062 21692 3068
rect 21548 2440 21600 2446
rect 21548 2382 21600 2388
rect 21088 2304 21140 2310
rect 21088 2246 21140 2252
rect 19350 2150 19354 2202
rect 19406 2150 19410 2202
rect 12716 1896 12768 1902
rect 12716 1838 12768 1844
rect 13268 1896 13320 1902
rect 13268 1838 13320 1844
rect 11612 1760 11664 1766
rect 11612 1702 11664 1708
rect 11350 1606 11354 1658
rect 11406 1606 11410 1658
rect 11350 1040 11410 1606
rect 11520 1556 11572 1562
rect 11440 1516 11520 1544
rect 11440 800 11468 1516
rect 11520 1498 11572 1504
rect 11624 800 11652 1702
rect 12164 1488 12216 1494
rect 12164 1430 12216 1436
rect 11980 1420 12032 1426
rect 11980 1362 12032 1368
rect 11992 800 12020 1362
rect 12176 800 12204 1430
rect 12348 1420 12400 1426
rect 12348 1362 12400 1368
rect 12360 800 12388 1362
rect 12728 800 12756 1838
rect 12900 1420 12952 1426
rect 12900 1362 12952 1368
rect 12912 800 12940 1362
rect 13280 800 13308 1838
rect 13452 1760 13504 1766
rect 13452 1702 13504 1708
rect 13820 1760 13872 1766
rect 13820 1702 13872 1708
rect 14556 1760 14608 1766
rect 14556 1702 14608 1708
rect 16948 1760 17000 1766
rect 16948 1702 17000 1708
rect 18236 1760 18288 1766
rect 18236 1702 18288 1708
rect 13464 800 13492 1702
rect 13832 800 13860 1702
rect 14004 1556 14056 1562
rect 14004 1498 14056 1504
rect 14016 800 14044 1498
rect 14188 1420 14240 1426
rect 14188 1362 14240 1368
rect 14200 800 14228 1362
rect 14568 800 14596 1702
rect 16212 1488 16264 1494
rect 16212 1430 16264 1436
rect 14740 1420 14792 1426
rect 14740 1362 14792 1368
rect 15108 1420 15160 1426
rect 15108 1362 15160 1368
rect 15292 1420 15344 1426
rect 15292 1362 15344 1368
rect 15660 1420 15712 1426
rect 15660 1362 15712 1368
rect 15844 1420 15896 1426
rect 15844 1362 15896 1368
rect 14752 800 14780 1362
rect 15120 800 15148 1362
rect 15304 800 15332 1362
rect 15672 800 15700 1362
rect 15856 800 15884 1362
rect 16224 800 16252 1430
rect 16396 1420 16448 1426
rect 16396 1362 16448 1368
rect 16580 1420 16632 1426
rect 16580 1362 16632 1368
rect 16408 800 16436 1362
rect 16592 800 16620 1362
rect 16960 800 16988 1702
rect 17684 1488 17736 1494
rect 17684 1430 17736 1436
rect 17132 1420 17184 1426
rect 17132 1362 17184 1368
rect 17500 1420 17552 1426
rect 17500 1362 17552 1368
rect 17144 800 17172 1362
rect 17512 800 17540 1362
rect 17696 800 17724 1430
rect 18144 1420 18196 1426
rect 18064 1380 18144 1408
rect 18064 800 18092 1380
rect 18144 1362 18196 1368
rect 18248 800 18276 1702
rect 18788 1556 18840 1562
rect 18788 1498 18840 1504
rect 18604 1488 18656 1494
rect 18604 1430 18656 1436
rect 18616 800 18644 1430
rect 18800 800 18828 1498
rect 18972 1420 19024 1426
rect 18972 1362 19024 1368
rect 18984 800 19012 1362
rect 19350 1268 19410 2150
rect 21100 1970 21128 2246
rect 21088 1964 21140 1970
rect 21088 1906 21140 1912
rect 20628 1896 20680 1902
rect 20628 1838 20680 1844
rect 19524 1760 19576 1766
rect 19524 1702 19576 1708
rect 20352 1760 20404 1766
rect 20352 1702 20404 1708
rect 19536 1578 19564 1702
rect 19350 1212 19352 1268
rect 19408 1212 19410 1268
rect 19350 1114 19410 1212
rect 19350 1062 19354 1114
rect 19406 1062 19410 1114
rect 19350 1040 19410 1062
rect 19444 1550 19564 1578
rect 20076 1556 20128 1562
rect 19444 898 19472 1550
rect 20076 1498 20128 1504
rect 19892 1488 19944 1494
rect 19892 1430 19944 1436
rect 19524 1420 19576 1426
rect 19524 1362 19576 1368
rect 19352 870 19472 898
rect 19352 800 19380 870
rect 19536 800 19564 1362
rect 19904 800 19932 1430
rect 20088 800 20116 1498
rect 20364 1426 20392 1702
rect 20352 1420 20404 1426
rect 20352 1362 20404 1368
rect 20444 1420 20496 1426
rect 20444 1362 20496 1368
rect 20456 800 20484 1362
rect 20640 800 20668 1838
rect 21180 1828 21232 1834
rect 21180 1770 21232 1776
rect 20996 1420 21048 1426
rect 20996 1362 21048 1368
rect 21008 800 21036 1362
rect 21192 800 21220 1770
rect 21652 1442 21680 3062
rect 21744 2650 21772 3800
rect 21732 2644 21784 2650
rect 21732 2586 21784 2592
rect 22112 1986 22140 3800
rect 22192 3392 22244 3398
rect 22192 3334 22244 3340
rect 22204 3058 22232 3334
rect 22192 3052 22244 3058
rect 22192 2994 22244 3000
rect 22296 2582 22324 3800
rect 22560 3460 22612 3466
rect 22560 3402 22612 3408
rect 22572 3058 22600 3402
rect 22560 3052 22612 3058
rect 22560 2994 22612 3000
rect 22468 2984 22520 2990
rect 22468 2926 22520 2932
rect 22284 2576 22336 2582
rect 22284 2518 22336 2524
rect 22020 1970 22140 1986
rect 22008 1964 22140 1970
rect 22060 1958 22140 1964
rect 22008 1906 22060 1912
rect 22008 1828 22060 1834
rect 22008 1770 22060 1776
rect 21732 1760 21784 1766
rect 21732 1702 21784 1708
rect 21376 1414 21680 1442
rect 21376 800 21404 1414
rect 21744 800 21772 1702
rect 22020 898 22048 1770
rect 22284 1488 22336 1494
rect 22284 1430 22336 1436
rect 21928 870 22048 898
rect 21928 800 21956 870
rect 22296 800 22324 1430
rect 22480 800 22508 2926
rect 22664 2650 22692 3800
rect 22652 2644 22704 2650
rect 22652 2586 22704 2592
rect 22848 1970 22876 3800
rect 23216 2514 23244 3800
rect 23400 2582 23428 3800
rect 23768 2650 23796 3800
rect 23952 2650 23980 3800
rect 23756 2644 23808 2650
rect 23756 2586 23808 2592
rect 23940 2644 23992 2650
rect 23940 2586 23992 2592
rect 24136 2582 24164 3800
rect 24504 3058 24532 3800
rect 24492 3052 24544 3058
rect 24492 2994 24544 3000
rect 23388 2576 23440 2582
rect 23388 2518 23440 2524
rect 24124 2576 24176 2582
rect 24124 2518 24176 2524
rect 24688 2514 24716 3800
rect 25056 2666 25084 3800
rect 24780 2650 25084 2666
rect 25240 2650 25268 3800
rect 25608 2650 25636 3800
rect 25792 3058 25820 3800
rect 25780 3052 25832 3058
rect 25780 2994 25832 3000
rect 25976 2938 26004 3800
rect 25792 2910 26004 2938
rect 25792 2650 25820 2910
rect 25872 2848 25924 2854
rect 25872 2790 25924 2796
rect 24768 2644 25084 2650
rect 24820 2638 25084 2644
rect 25228 2644 25280 2650
rect 24768 2586 24820 2592
rect 25228 2586 25280 2592
rect 25596 2644 25648 2650
rect 25596 2586 25648 2592
rect 25780 2644 25832 2650
rect 25780 2586 25832 2592
rect 25502 2544 25558 2553
rect 23204 2508 23256 2514
rect 23204 2450 23256 2456
rect 24676 2508 24728 2514
rect 24676 2450 24728 2456
rect 24768 2508 24820 2514
rect 25502 2479 25558 2488
rect 24768 2450 24820 2456
rect 22928 2440 22980 2446
rect 22928 2382 22980 2388
rect 22836 1964 22888 1970
rect 22836 1906 22888 1912
rect 22836 1828 22888 1834
rect 22836 1770 22888 1776
rect 22848 800 22876 1770
rect 22940 1562 22968 2382
rect 23112 2372 23164 2378
rect 23112 2314 23164 2320
rect 23124 1970 23152 2314
rect 23848 2100 23900 2106
rect 23848 2042 23900 2048
rect 23296 2032 23348 2038
rect 23294 2000 23296 2009
rect 23348 2000 23350 2009
rect 23112 1964 23164 1970
rect 23294 1935 23350 1944
rect 23112 1906 23164 1912
rect 23572 1828 23624 1834
rect 23572 1770 23624 1776
rect 22928 1556 22980 1562
rect 22928 1498 22980 1504
rect 23020 1556 23072 1562
rect 23020 1498 23072 1504
rect 23032 800 23060 1498
rect 23388 1352 23440 1358
rect 23388 1294 23440 1300
rect 23400 800 23428 1294
rect 23584 800 23612 1770
rect 23756 1488 23808 1494
rect 23756 1430 23808 1436
rect 23768 800 23796 1430
rect 23860 1358 23888 2042
rect 24780 1970 24808 2450
rect 25516 2446 25544 2479
rect 25504 2440 25556 2446
rect 25504 2382 25556 2388
rect 25596 2440 25648 2446
rect 25596 2382 25648 2388
rect 25044 2372 25096 2378
rect 25044 2314 25096 2320
rect 24952 2304 25004 2310
rect 24952 2246 25004 2252
rect 24768 1964 24820 1970
rect 24768 1906 24820 1912
rect 24400 1896 24452 1902
rect 24136 1844 24400 1850
rect 24136 1838 24452 1844
rect 24136 1822 24440 1838
rect 23848 1352 23900 1358
rect 23848 1294 23900 1300
rect 24136 800 24164 1822
rect 24308 1760 24360 1766
rect 24308 1702 24360 1708
rect 24320 800 24348 1702
rect 24768 1488 24820 1494
rect 24688 1448 24768 1476
rect 24688 800 24716 1448
rect 24768 1430 24820 1436
rect 24964 898 24992 2246
rect 25056 1970 25084 2314
rect 25320 2304 25372 2310
rect 25320 2246 25372 2252
rect 25226 2000 25282 2009
rect 25044 1964 25096 1970
rect 25332 1970 25360 2246
rect 25608 1970 25636 2382
rect 25226 1935 25282 1944
rect 25320 1964 25372 1970
rect 25044 1906 25096 1912
rect 25042 1592 25098 1601
rect 25042 1527 25044 1536
rect 25096 1527 25098 1536
rect 25044 1498 25096 1504
rect 24872 870 24992 898
rect 24872 800 24900 870
rect 25240 800 25268 1935
rect 25320 1906 25372 1912
rect 25596 1964 25648 1970
rect 25596 1906 25648 1912
rect 25884 1442 25912 2790
rect 26344 2650 26372 3800
rect 26528 2650 26556 3800
rect 26332 2644 26384 2650
rect 26332 2586 26384 2592
rect 26516 2644 26568 2650
rect 26516 2586 26568 2592
rect 26896 2582 26924 3800
rect 27080 2650 27108 3800
rect 27350 2746 27410 3312
rect 27350 2694 27354 2746
rect 27406 2694 27410 2746
rect 27068 2644 27120 2650
rect 27068 2586 27120 2592
rect 26056 2576 26108 2582
rect 26148 2576 26200 2582
rect 26056 2518 26108 2524
rect 26146 2544 26148 2553
rect 26424 2576 26476 2582
rect 26200 2544 26202 2553
rect 25964 1760 26016 1766
rect 25964 1702 26016 1708
rect 25976 1601 26004 1702
rect 25962 1592 26018 1601
rect 25962 1527 26018 1536
rect 25884 1414 26004 1442
rect 25780 1284 25832 1290
rect 25780 1226 25832 1232
rect 25412 1216 25464 1222
rect 25412 1158 25464 1164
rect 25424 800 25452 1158
rect 25792 800 25820 1226
rect 25976 800 26004 1414
rect 26068 898 26096 2518
rect 26884 2576 26936 2582
rect 26476 2524 26556 2530
rect 26424 2518 26556 2524
rect 26884 2518 26936 2524
rect 26146 2479 26202 2488
rect 26240 2508 26292 2514
rect 26436 2502 26556 2518
rect 26240 2450 26292 2456
rect 26148 2032 26200 2038
rect 26148 1974 26200 1980
rect 26160 1222 26188 1974
rect 26252 1834 26280 2450
rect 26332 2032 26384 2038
rect 26332 1974 26384 1980
rect 26240 1828 26292 1834
rect 26240 1770 26292 1776
rect 26344 1494 26372 1974
rect 26332 1488 26384 1494
rect 26332 1430 26384 1436
rect 26148 1216 26200 1222
rect 26148 1158 26200 1164
rect 26068 870 26188 898
rect 26160 800 26188 870
rect 26528 800 26556 2502
rect 27350 2348 27410 2694
rect 27448 2564 27476 3800
rect 27632 2650 27660 3800
rect 28000 3058 28028 3800
rect 27988 3052 28040 3058
rect 27988 2994 28040 3000
rect 28184 2650 28212 3800
rect 27620 2644 27672 2650
rect 27620 2586 27672 2592
rect 28172 2644 28224 2650
rect 28172 2586 28224 2592
rect 27528 2576 27580 2582
rect 27448 2536 27528 2564
rect 27528 2518 27580 2524
rect 28264 2508 28316 2514
rect 28264 2450 28316 2456
rect 27350 2292 27352 2348
rect 27408 2292 27410 2348
rect 27804 2372 27856 2378
rect 27804 2314 27856 2320
rect 27068 2100 27120 2106
rect 27068 2042 27120 2048
rect 26608 1964 26660 1970
rect 26608 1906 26660 1912
rect 26620 1494 26648 1906
rect 26608 1488 26660 1494
rect 26608 1430 26660 1436
rect 26700 1216 26752 1222
rect 26700 1158 26752 1164
rect 26712 800 26740 1158
rect 27080 800 27108 2042
rect 27252 1828 27304 1834
rect 27252 1770 27304 1776
rect 27264 800 27292 1770
rect 27350 1658 27410 2292
rect 27712 2032 27764 2038
rect 27712 1974 27764 1980
rect 27350 1606 27354 1658
rect 27406 1606 27410 1658
rect 27350 1040 27410 1606
rect 27724 1562 27752 1974
rect 27620 1556 27672 1562
rect 27620 1498 27672 1504
rect 27712 1556 27764 1562
rect 27712 1498 27764 1504
rect 27632 800 27660 1498
rect 27816 800 27844 2314
rect 27896 1760 27948 1766
rect 27948 1720 28028 1748
rect 27896 1702 27948 1708
rect 28000 800 28028 1720
rect 28276 1442 28304 2450
rect 28368 2446 28396 3800
rect 28736 3058 28764 3800
rect 28724 3052 28776 3058
rect 28724 2994 28776 3000
rect 28920 2582 28948 3800
rect 29288 2922 29316 3800
rect 29276 2916 29328 2922
rect 29276 2858 29328 2864
rect 29472 2650 29500 3800
rect 29460 2644 29512 2650
rect 29460 2586 29512 2592
rect 29840 2582 29868 3800
rect 30024 2650 30052 3800
rect 30392 2650 30420 3800
rect 30012 2644 30064 2650
rect 30012 2586 30064 2592
rect 30380 2644 30432 2650
rect 30380 2586 30432 2592
rect 30576 2582 30604 3800
rect 30760 2650 30788 3800
rect 30748 2644 30800 2650
rect 30748 2586 30800 2592
rect 28908 2576 28960 2582
rect 28908 2518 28960 2524
rect 29828 2576 29880 2582
rect 29828 2518 29880 2524
rect 30564 2576 30616 2582
rect 30564 2518 30616 2524
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 28448 2372 28500 2378
rect 28448 2314 28500 2320
rect 28460 1562 28488 2314
rect 28540 2304 28592 2310
rect 28540 2246 28592 2252
rect 30380 2304 30432 2310
rect 30380 2246 30432 2252
rect 28448 1556 28500 1562
rect 28448 1498 28500 1504
rect 28276 1414 28396 1442
rect 28368 800 28396 1414
rect 28552 800 28580 2246
rect 29460 2100 29512 2106
rect 29460 2042 29512 2048
rect 29552 2100 29604 2106
rect 29552 2042 29604 2048
rect 28816 1828 28868 1834
rect 28816 1770 28868 1776
rect 28828 1714 28856 1770
rect 29092 1760 29144 1766
rect 28828 1686 29040 1714
rect 29092 1702 29144 1708
rect 28816 1284 28868 1290
rect 28868 1244 28948 1272
rect 28816 1226 28868 1232
rect 28920 800 28948 1244
rect 29012 898 29040 1686
rect 29104 1562 29132 1702
rect 29092 1556 29144 1562
rect 29092 1498 29144 1504
rect 29012 870 29132 898
rect 29104 800 29132 870
rect 29472 800 29500 2042
rect 29564 1358 29592 2042
rect 30392 1970 30420 2246
rect 30656 2032 30708 2038
rect 30656 1974 30708 1980
rect 30932 2032 30984 2038
rect 30932 1974 30984 1980
rect 29644 1964 29696 1970
rect 29644 1906 29696 1912
rect 30380 1964 30432 1970
rect 30380 1906 30432 1912
rect 29552 1352 29604 1358
rect 29552 1294 29604 1300
rect 29656 800 29684 1906
rect 30012 1760 30064 1766
rect 30012 1702 30064 1708
rect 30564 1760 30616 1766
rect 30564 1702 30616 1708
rect 30024 800 30052 1702
rect 30576 1562 30604 1702
rect 30564 1556 30616 1562
rect 30564 1498 30616 1504
rect 30196 1420 30248 1426
rect 30196 1362 30248 1368
rect 30208 800 30236 1362
rect 30380 1216 30432 1222
rect 30380 1158 30432 1164
rect 30392 800 30420 1158
rect 30668 898 30696 1974
rect 30840 1896 30892 1902
rect 30840 1838 30892 1844
rect 30748 1828 30800 1834
rect 30748 1770 30800 1776
rect 30760 1494 30788 1770
rect 30748 1488 30800 1494
rect 30748 1430 30800 1436
rect 30852 898 30880 1838
rect 30944 1494 30972 1974
rect 31128 1970 31156 3800
rect 31312 2650 31340 3800
rect 31576 3596 31628 3602
rect 31576 3538 31628 3544
rect 31588 3058 31616 3538
rect 31576 3052 31628 3058
rect 31576 2994 31628 3000
rect 31300 2644 31352 2650
rect 31300 2586 31352 2592
rect 31680 2582 31708 3800
rect 31668 2576 31720 2582
rect 31668 2518 31720 2524
rect 31864 2446 31892 3800
rect 32232 2514 32260 3800
rect 32416 2922 32444 3800
rect 32784 3058 32812 3800
rect 32772 3052 32824 3058
rect 32772 2994 32824 3000
rect 32404 2916 32456 2922
rect 32404 2858 32456 2864
rect 32968 2582 32996 3800
rect 33048 2644 33100 2650
rect 33152 2632 33180 3800
rect 33232 3528 33284 3534
rect 33232 3470 33284 3476
rect 33244 3058 33272 3470
rect 33232 3052 33284 3058
rect 33232 2994 33284 3000
rect 33520 2650 33548 3800
rect 33100 2604 33180 2632
rect 33508 2644 33560 2650
rect 33048 2586 33100 2592
rect 33508 2586 33560 2592
rect 33704 2582 33732 3800
rect 33784 3460 33836 3466
rect 33784 3402 33836 3408
rect 33796 3058 33824 3402
rect 33784 3052 33836 3058
rect 33784 2994 33836 3000
rect 32956 2576 33008 2582
rect 32956 2518 33008 2524
rect 33692 2576 33744 2582
rect 33692 2518 33744 2524
rect 34072 2514 34100 3800
rect 34256 2650 34284 3800
rect 34624 3482 34652 3800
rect 34348 3454 34652 3482
rect 34348 3194 34376 3454
rect 34520 3392 34572 3398
rect 34520 3334 34572 3340
rect 34532 3210 34560 3334
rect 34336 3188 34388 3194
rect 34336 3130 34388 3136
rect 34440 3182 34560 3210
rect 34440 3126 34468 3182
rect 34428 3120 34480 3126
rect 34428 3062 34480 3068
rect 34808 2854 34836 3800
rect 35176 3602 35204 3800
rect 35164 3596 35216 3602
rect 35164 3538 35216 3544
rect 35360 3448 35388 3800
rect 35176 3420 35388 3448
rect 35176 2990 35204 3420
rect 35544 3398 35572 3800
rect 35912 3534 35940 3800
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 36096 3466 36124 3800
rect 36084 3460 36136 3466
rect 36084 3402 36136 3408
rect 36176 3460 36228 3466
rect 36176 3402 36228 3408
rect 35532 3392 35584 3398
rect 35532 3334 35584 3340
rect 35350 3290 35410 3312
rect 35350 3238 35354 3290
rect 35406 3238 35410 3290
rect 35164 2984 35216 2990
rect 35164 2926 35216 2932
rect 34796 2848 34848 2854
rect 34796 2790 34848 2796
rect 34244 2644 34296 2650
rect 34244 2586 34296 2592
rect 32220 2508 32272 2514
rect 32220 2450 32272 2456
rect 34060 2508 34112 2514
rect 34060 2450 34112 2456
rect 31852 2440 31904 2446
rect 31852 2382 31904 2388
rect 31300 2372 31352 2378
rect 31300 2314 31352 2320
rect 31116 1964 31168 1970
rect 31116 1906 31168 1912
rect 30932 1488 30984 1494
rect 30932 1430 30984 1436
rect 30668 870 30788 898
rect 30852 870 30972 898
rect 30760 800 30788 870
rect 30944 800 30972 870
rect 31312 800 31340 2314
rect 33140 2304 33192 2310
rect 33140 2246 33192 2252
rect 32404 2100 32456 2106
rect 32404 2042 32456 2048
rect 31392 1964 31444 1970
rect 31392 1906 31444 1912
rect 31404 1562 31432 1906
rect 31576 1896 31628 1902
rect 31576 1838 31628 1844
rect 31484 1828 31536 1834
rect 31484 1770 31536 1776
rect 31392 1556 31444 1562
rect 31392 1498 31444 1504
rect 31496 800 31524 1770
rect 31588 1562 31616 1838
rect 31760 1828 31812 1834
rect 31760 1770 31812 1776
rect 32220 1828 32272 1834
rect 32220 1770 32272 1776
rect 31576 1556 31628 1562
rect 31576 1498 31628 1504
rect 31772 1358 31800 1770
rect 32036 1760 32088 1766
rect 32036 1702 32088 1708
rect 31760 1352 31812 1358
rect 31760 1294 31812 1300
rect 31760 1216 31812 1222
rect 31812 1176 31892 1204
rect 31760 1158 31812 1164
rect 31864 800 31892 1176
rect 32048 800 32076 1702
rect 32232 1562 32260 1770
rect 32220 1556 32272 1562
rect 32220 1498 32272 1504
rect 32416 800 32444 2042
rect 32772 1760 32824 1766
rect 32772 1702 32824 1708
rect 32864 1760 32916 1766
rect 32864 1702 32916 1708
rect 32588 1420 32640 1426
rect 32588 1362 32640 1368
rect 32600 800 32628 1362
rect 32784 800 32812 1702
rect 32876 1426 32904 1702
rect 32864 1420 32916 1426
rect 32864 1362 32916 1368
rect 33152 800 33180 2246
rect 35350 2202 35410 3238
rect 35728 2922 35848 2938
rect 35728 2916 35860 2922
rect 35728 2910 35808 2916
rect 35624 2848 35676 2854
rect 35728 2836 35756 2910
rect 35808 2858 35860 2864
rect 36188 2854 36216 3402
rect 36464 2922 36492 3800
rect 36648 3194 36676 3800
rect 37016 3466 37044 3800
rect 37004 3460 37056 3466
rect 37004 3402 37056 3408
rect 36912 3392 36964 3398
rect 36912 3334 36964 3340
rect 36636 3188 36688 3194
rect 36636 3130 36688 3136
rect 36924 2922 36952 3334
rect 37200 2990 37228 3800
rect 37280 3460 37332 3466
rect 37280 3402 37332 3408
rect 37188 2984 37240 2990
rect 37188 2926 37240 2932
rect 36452 2916 36504 2922
rect 36452 2858 36504 2864
rect 36912 2916 36964 2922
rect 36912 2858 36964 2864
rect 35676 2808 35756 2836
rect 36176 2848 36228 2854
rect 35624 2790 35676 2796
rect 36176 2790 36228 2796
rect 37096 2848 37148 2854
rect 37292 2802 37320 3402
rect 37568 3058 37596 3800
rect 37752 3126 37780 3800
rect 37740 3120 37792 3126
rect 37740 3062 37792 3068
rect 37556 3052 37608 3058
rect 37556 2994 37608 3000
rect 37148 2796 37320 2802
rect 37096 2790 37320 2796
rect 37108 2774 37320 2790
rect 37936 2650 37964 3800
rect 38304 3466 38332 3800
rect 38292 3460 38344 3466
rect 38292 3402 38344 3408
rect 38488 3194 38516 3800
rect 38856 3618 38884 3800
rect 38764 3590 38884 3618
rect 38764 3398 38792 3590
rect 38844 3460 38896 3466
rect 38844 3402 38896 3408
rect 38752 3392 38804 3398
rect 38752 3334 38804 3340
rect 38476 3188 38528 3194
rect 38476 3130 38528 3136
rect 38660 3188 38712 3194
rect 38660 3130 38712 3136
rect 38672 2854 38700 3130
rect 38856 2854 38884 3402
rect 39040 3126 39068 3800
rect 39120 3392 39172 3398
rect 39120 3334 39172 3340
rect 39028 3120 39080 3126
rect 39028 3062 39080 3068
rect 39132 2854 39160 3334
rect 39408 3058 39436 3800
rect 39592 3194 39620 3800
rect 39580 3188 39632 3194
rect 39580 3130 39632 3136
rect 39396 3052 39448 3058
rect 39396 2994 39448 3000
rect 39488 3052 39540 3058
rect 39488 2994 39540 3000
rect 39500 2854 39528 2994
rect 39776 2922 39804 3800
rect 40144 2990 40172 3800
rect 40132 2984 40184 2990
rect 40132 2926 40184 2932
rect 39764 2916 39816 2922
rect 39764 2858 39816 2864
rect 38660 2848 38712 2854
rect 38660 2790 38712 2796
rect 38844 2848 38896 2854
rect 38844 2790 38896 2796
rect 39120 2848 39172 2854
rect 39120 2790 39172 2796
rect 39488 2848 39540 2854
rect 39488 2790 39540 2796
rect 40328 2650 40356 3800
rect 40696 3466 40724 3800
rect 40684 3460 40736 3466
rect 40684 3402 40736 3408
rect 40880 3398 40908 3800
rect 40868 3392 40920 3398
rect 40868 3334 40920 3340
rect 41248 2990 41276 3800
rect 41236 2984 41288 2990
rect 41236 2926 41288 2932
rect 41432 2854 41460 3800
rect 41800 2922 41828 3800
rect 41984 3058 42012 3800
rect 42168 3194 42196 3800
rect 42156 3188 42208 3194
rect 42156 3130 42208 3136
rect 42536 3126 42564 3800
rect 42524 3120 42576 3126
rect 42524 3062 42576 3068
rect 41972 3052 42024 3058
rect 41972 2994 42024 3000
rect 41788 2916 41840 2922
rect 41788 2858 41840 2864
rect 41420 2848 41472 2854
rect 41420 2790 41472 2796
rect 37924 2644 37976 2650
rect 37924 2586 37976 2592
rect 40316 2644 40368 2650
rect 40316 2586 40368 2592
rect 42720 2582 42748 3800
rect 42800 3392 42852 3398
rect 42800 3334 42852 3340
rect 42812 3058 42840 3334
rect 42800 3052 42852 3058
rect 42800 2994 42852 3000
rect 43088 2990 43116 3800
rect 43272 3398 43300 3800
rect 43260 3392 43312 3398
rect 43260 3334 43312 3340
rect 43076 2984 43128 2990
rect 43076 2926 43128 2932
rect 43350 2746 43410 3312
rect 43350 2694 43354 2746
rect 43406 2694 43410 2746
rect 42708 2576 42760 2582
rect 42708 2518 42760 2524
rect 35350 2150 35354 2202
rect 35406 2150 35410 2202
rect 33692 2032 33744 2038
rect 33692 1974 33744 1980
rect 34152 2032 34204 2038
rect 34152 1974 34204 1980
rect 33324 1964 33376 1970
rect 33324 1906 33376 1912
rect 33336 800 33364 1906
rect 33704 800 33732 1974
rect 34164 1562 34192 1974
rect 34796 1964 34848 1970
rect 34796 1906 34848 1912
rect 34244 1896 34296 1902
rect 34244 1838 34296 1844
rect 34428 1896 34480 1902
rect 34428 1838 34480 1844
rect 33784 1556 33836 1562
rect 33784 1498 33836 1504
rect 34152 1556 34204 1562
rect 34152 1498 34204 1504
rect 33796 898 33824 1498
rect 33796 870 33916 898
rect 33888 800 33916 870
rect 34256 800 34284 1838
rect 34440 1562 34468 1838
rect 34704 1828 34756 1834
rect 34704 1770 34756 1776
rect 34428 1556 34480 1562
rect 34428 1498 34480 1504
rect 34428 1216 34480 1222
rect 34428 1158 34480 1164
rect 34440 800 34468 1158
rect 34716 898 34744 1770
rect 34808 1562 34836 1906
rect 35072 1828 35124 1834
rect 35072 1770 35124 1776
rect 35084 1562 35112 1770
rect 35164 1760 35216 1766
rect 35164 1702 35216 1708
rect 34796 1556 34848 1562
rect 34796 1498 34848 1504
rect 35072 1556 35124 1562
rect 35072 1498 35124 1504
rect 34980 1352 35032 1358
rect 34980 1294 35032 1300
rect 34716 870 34836 898
rect 34808 800 34836 870
rect 34992 800 35020 1294
rect 35176 800 35204 1702
rect 35350 1268 35410 2150
rect 43350 2348 43410 2694
rect 43640 2650 43668 3800
rect 43824 2922 43852 3800
rect 43812 2916 43864 2922
rect 43812 2858 43864 2864
rect 44192 2854 44220 3800
rect 44272 3392 44324 3398
rect 44272 3334 44324 3340
rect 44284 3058 44312 3334
rect 44376 3194 44404 3800
rect 44364 3188 44416 3194
rect 44364 3130 44416 3136
rect 44560 3126 44588 3800
rect 44548 3120 44600 3126
rect 44548 3062 44600 3068
rect 44272 3052 44324 3058
rect 44272 2994 44324 3000
rect 44928 2922 44956 3800
rect 45112 3398 45140 3800
rect 45100 3392 45152 3398
rect 45100 3334 45152 3340
rect 44916 2916 44968 2922
rect 44916 2858 44968 2864
rect 45480 2854 45508 3800
rect 45664 2990 45692 3800
rect 45652 2984 45704 2990
rect 45652 2926 45704 2932
rect 44180 2848 44232 2854
rect 44180 2790 44232 2796
rect 45468 2848 45520 2854
rect 45468 2790 45520 2796
rect 43628 2644 43680 2650
rect 43628 2586 43680 2592
rect 46032 2582 46060 3800
rect 46216 3194 46244 3800
rect 46204 3188 46256 3194
rect 46204 3130 46256 3136
rect 46584 2650 46612 3800
rect 46768 3058 46796 3800
rect 46952 3126 46980 3800
rect 46940 3120 46992 3126
rect 46940 3062 46992 3068
rect 46756 3052 46808 3058
rect 46756 2994 46808 3000
rect 47216 2848 47268 2854
rect 47320 2836 47348 3800
rect 47504 2990 47532 3800
rect 47492 2984 47544 2990
rect 47492 2926 47544 2932
rect 47872 2922 47900 3800
rect 48056 3058 48084 3800
rect 48044 3052 48096 3058
rect 48044 2994 48096 3000
rect 47860 2916 47912 2922
rect 47860 2858 47912 2864
rect 47268 2808 47348 2836
rect 47216 2790 47268 2796
rect 48424 2666 48452 3800
rect 48608 3126 48636 3800
rect 48596 3120 48648 3126
rect 48596 3062 48648 3068
rect 48976 3058 49004 3800
rect 48964 3052 49016 3058
rect 48964 2994 49016 3000
rect 48240 2650 48452 2666
rect 46572 2644 46624 2650
rect 46572 2586 46624 2592
rect 48228 2644 48452 2650
rect 48280 2638 48452 2644
rect 48228 2586 48280 2592
rect 49160 2582 49188 3800
rect 49344 2854 49372 3800
rect 49712 2922 49740 3800
rect 49896 2990 49924 3800
rect 50264 3058 50292 3800
rect 50448 3126 50476 3800
rect 50436 3120 50488 3126
rect 50436 3062 50488 3068
rect 50252 3052 50304 3058
rect 50252 2994 50304 3000
rect 50816 2990 50844 3800
rect 49884 2984 49936 2990
rect 49884 2926 49936 2932
rect 50804 2984 50856 2990
rect 50804 2926 50856 2932
rect 51000 2922 51028 3800
rect 51368 3380 51396 3800
rect 51092 3352 51396 3380
rect 49700 2916 49752 2922
rect 49700 2858 49752 2864
rect 50988 2916 51040 2922
rect 50988 2858 51040 2864
rect 49332 2848 49384 2854
rect 49332 2790 49384 2796
rect 51092 2666 51120 3352
rect 51000 2650 51120 2666
rect 50988 2644 51120 2650
rect 51040 2638 51120 2644
rect 51350 3290 51410 3312
rect 51350 3238 51354 3290
rect 51406 3238 51410 3290
rect 50988 2586 51040 2592
rect 46020 2576 46072 2582
rect 46020 2518 46072 2524
rect 49148 2576 49200 2582
rect 49148 2518 49200 2524
rect 43350 2292 43352 2348
rect 43408 2292 43410 2348
rect 36268 2100 36320 2106
rect 36268 2042 36320 2048
rect 35716 1760 35768 1766
rect 35716 1702 35768 1708
rect 35728 1562 35756 1702
rect 35532 1556 35584 1562
rect 35532 1498 35584 1504
rect 35716 1556 35768 1562
rect 35716 1498 35768 1504
rect 35350 1212 35352 1268
rect 35408 1212 35410 1268
rect 35350 1114 35410 1212
rect 35350 1062 35354 1114
rect 35406 1062 35410 1114
rect 35350 1040 35410 1062
rect 35544 800 35572 1498
rect 35716 1284 35768 1290
rect 35716 1226 35768 1232
rect 35728 800 35756 1226
rect 36084 1216 36136 1222
rect 36084 1158 36136 1164
rect 36096 800 36124 1158
rect 36280 800 36308 2042
rect 36636 2032 36688 2038
rect 36636 1974 36688 1980
rect 38200 2032 38252 2038
rect 38200 1974 38252 1980
rect 40132 2032 40184 2038
rect 40132 1974 40184 1980
rect 36648 800 36676 1974
rect 37188 1964 37240 1970
rect 37188 1906 37240 1912
rect 36820 1896 36872 1902
rect 36820 1838 36872 1844
rect 36832 800 36860 1838
rect 37200 800 37228 1906
rect 37280 1896 37332 1902
rect 37280 1838 37332 1844
rect 37292 1562 37320 1838
rect 37372 1828 37424 1834
rect 37372 1770 37424 1776
rect 37648 1828 37700 1834
rect 37648 1770 37700 1776
rect 37280 1556 37332 1562
rect 37280 1498 37332 1504
rect 37384 800 37412 1770
rect 37660 1494 37688 1770
rect 37832 1760 37884 1766
rect 37884 1720 37964 1748
rect 37832 1702 37884 1708
rect 37556 1488 37608 1494
rect 37556 1430 37608 1436
rect 37648 1488 37700 1494
rect 37648 1430 37700 1436
rect 37568 800 37596 1430
rect 37936 800 37964 1720
rect 38212 1358 38240 1974
rect 39028 1896 39080 1902
rect 39028 1838 39080 1844
rect 39672 1896 39724 1902
rect 39672 1838 39724 1844
rect 38476 1420 38528 1426
rect 38476 1362 38528 1368
rect 38108 1352 38160 1358
rect 38108 1294 38160 1300
rect 38200 1352 38252 1358
rect 38200 1294 38252 1300
rect 38120 800 38148 1294
rect 38488 800 38516 1362
rect 38660 1284 38712 1290
rect 38660 1226 38712 1232
rect 38672 800 38700 1226
rect 39040 800 39068 1838
rect 39120 1556 39172 1562
rect 39172 1516 39252 1544
rect 39120 1498 39172 1504
rect 39224 800 39252 1516
rect 39580 1488 39632 1494
rect 39580 1430 39632 1436
rect 39592 800 39620 1430
rect 39684 1358 39712 1838
rect 39764 1828 39816 1834
rect 39764 1770 39816 1776
rect 39672 1352 39724 1358
rect 39672 1294 39724 1300
rect 39776 800 39804 1770
rect 39948 1760 40000 1766
rect 39948 1702 40000 1708
rect 39960 800 39988 1702
rect 40144 898 40172 1974
rect 41420 1964 41472 1970
rect 41420 1906 41472 1912
rect 42064 1964 42116 1970
rect 42064 1906 42116 1912
rect 42708 1964 42760 1970
rect 42708 1906 42760 1912
rect 40224 1828 40276 1834
rect 40224 1770 40276 1776
rect 40236 1494 40264 1770
rect 41052 1556 41104 1562
rect 41052 1498 41104 1504
rect 40224 1488 40276 1494
rect 40224 1430 40276 1436
rect 40316 1352 40368 1358
rect 40316 1294 40368 1300
rect 40328 1170 40356 1294
rect 40868 1216 40920 1222
rect 40328 1142 40540 1170
rect 40868 1158 40920 1164
rect 40144 870 40356 898
rect 40328 800 40356 870
rect 40512 800 40540 1142
rect 40880 800 40908 1158
rect 41064 800 41092 1498
rect 41432 800 41460 1906
rect 41604 1896 41656 1902
rect 41604 1838 41656 1844
rect 41616 800 41644 1838
rect 42076 1494 42104 1906
rect 42156 1828 42208 1834
rect 42156 1770 42208 1776
rect 42064 1488 42116 1494
rect 42064 1430 42116 1436
rect 41788 1284 41840 1290
rect 41788 1226 41840 1232
rect 41800 800 41828 1226
rect 42168 800 42196 1770
rect 42340 1352 42392 1358
rect 42340 1294 42392 1300
rect 42352 800 42380 1294
rect 42720 800 42748 1906
rect 42892 1828 42944 1834
rect 42892 1770 42944 1776
rect 42800 1760 42852 1766
rect 42800 1702 42852 1708
rect 42812 898 42840 1702
rect 42904 1494 42932 1770
rect 43350 1658 43410 2292
rect 51350 2202 51410 3238
rect 51552 3058 51580 3800
rect 51736 3126 51764 3800
rect 51724 3120 51776 3126
rect 51724 3062 51776 3068
rect 51540 3052 51592 3058
rect 51540 2994 51592 3000
rect 52104 2650 52132 3800
rect 52288 2922 52316 3800
rect 52656 2990 52684 3800
rect 52840 3126 52868 3800
rect 52828 3120 52880 3126
rect 52828 3062 52880 3068
rect 52644 2984 52696 2990
rect 52644 2926 52696 2932
rect 53208 2922 53236 3800
rect 53392 2990 53420 3800
rect 53576 3058 53604 3800
rect 53564 3052 53616 3058
rect 53564 2994 53616 3000
rect 53380 2984 53432 2990
rect 53380 2926 53432 2932
rect 52276 2916 52328 2922
rect 52276 2858 52328 2864
rect 53196 2916 53248 2922
rect 53196 2858 53248 2864
rect 53944 2666 53972 3800
rect 54128 2922 54156 3800
rect 54496 3126 54524 3800
rect 54484 3120 54536 3126
rect 54484 3062 54536 3068
rect 54680 3058 54708 3800
rect 54668 3052 54720 3058
rect 54668 2994 54720 3000
rect 55048 2922 55076 3800
rect 55232 2990 55260 3800
rect 55600 3058 55628 3800
rect 55588 3052 55640 3058
rect 55588 2994 55640 3000
rect 55220 2984 55272 2990
rect 55220 2926 55272 2932
rect 54116 2916 54168 2922
rect 54116 2858 54168 2864
rect 55036 2916 55088 2922
rect 55036 2858 55088 2864
rect 55678 2816 55734 2825
rect 55678 2751 55734 2760
rect 53760 2650 53972 2666
rect 52092 2644 52144 2650
rect 52092 2586 52144 2592
rect 53748 2644 53972 2650
rect 53800 2638 53972 2644
rect 53748 2586 53800 2592
rect 51350 2150 51354 2202
rect 51406 2150 51410 2202
rect 43996 1896 44048 1902
rect 43996 1838 44048 1844
rect 43812 1828 43864 1834
rect 43812 1770 43864 1776
rect 43350 1606 43354 1658
rect 43406 1606 43410 1658
rect 42892 1488 42944 1494
rect 42892 1430 42944 1436
rect 43260 1352 43312 1358
rect 43260 1294 43312 1300
rect 42812 870 42932 898
rect 42904 800 42932 870
rect 43272 800 43300 1294
rect 43350 1040 43410 1606
rect 43444 1556 43496 1562
rect 43444 1498 43496 1504
rect 43456 800 43484 1498
rect 43824 800 43852 1770
rect 44008 800 44036 1838
rect 46572 1828 46624 1834
rect 46572 1770 46624 1776
rect 44732 1760 44784 1766
rect 44732 1702 44784 1708
rect 45468 1760 45520 1766
rect 45468 1702 45520 1708
rect 44548 1488 44600 1494
rect 44548 1430 44600 1436
rect 44180 1420 44232 1426
rect 44180 1362 44232 1368
rect 44192 800 44220 1362
rect 44560 800 44588 1430
rect 44744 800 44772 1702
rect 45100 1488 45152 1494
rect 45100 1430 45152 1436
rect 45008 1216 45060 1222
rect 45008 1158 45060 1164
rect 45112 1170 45140 1430
rect 45480 1358 45508 1702
rect 46388 1556 46440 1562
rect 46388 1498 46440 1504
rect 46204 1488 46256 1494
rect 46204 1430 46256 1436
rect 45652 1420 45704 1426
rect 45652 1362 45704 1368
rect 45468 1352 45520 1358
rect 45468 1294 45520 1300
rect 45020 898 45048 1158
rect 45112 1142 45324 1170
rect 45020 870 45140 898
rect 45112 800 45140 870
rect 45296 800 45324 1142
rect 45664 800 45692 1362
rect 45836 1284 45888 1290
rect 45836 1226 45888 1232
rect 45848 800 45876 1226
rect 46216 800 46244 1430
rect 46400 800 46428 1498
rect 46584 800 46612 1770
rect 46940 1760 46992 1766
rect 46940 1702 46992 1708
rect 49516 1760 49568 1766
rect 49516 1702 49568 1708
rect 50988 1760 51040 1766
rect 50988 1702 51040 1708
rect 46952 800 46980 1702
rect 48044 1556 48096 1562
rect 48044 1498 48096 1504
rect 49240 1556 49292 1562
rect 49240 1498 49292 1504
rect 47032 1488 47084 1494
rect 47084 1448 47164 1476
rect 47032 1430 47084 1436
rect 47136 800 47164 1448
rect 47676 1420 47728 1426
rect 47676 1362 47728 1368
rect 47400 1352 47452 1358
rect 47452 1312 47532 1340
rect 47400 1294 47452 1300
rect 47504 800 47532 1312
rect 47688 800 47716 1362
rect 48056 800 48084 1498
rect 48228 1488 48280 1494
rect 48228 1430 48280 1436
rect 48964 1488 49016 1494
rect 48964 1430 49016 1436
rect 48240 800 48268 1430
rect 48596 1420 48648 1426
rect 48596 1362 48648 1368
rect 48608 800 48636 1362
rect 48780 1352 48832 1358
rect 48780 1294 48832 1300
rect 48792 800 48820 1294
rect 48976 800 49004 1430
rect 49252 898 49280 1498
rect 49252 870 49372 898
rect 49344 800 49372 870
rect 49528 800 49556 1702
rect 49988 1562 50476 1578
rect 49976 1556 50476 1562
rect 50028 1550 50476 1556
rect 49976 1498 50028 1504
rect 50068 1488 50120 1494
rect 50068 1430 50120 1436
rect 49884 1284 49936 1290
rect 49884 1226 49936 1232
rect 49896 800 49924 1226
rect 50080 800 50108 1430
rect 50448 800 50476 1550
rect 50620 1420 50672 1426
rect 50620 1362 50672 1368
rect 50632 800 50660 1362
rect 51000 800 51028 1702
rect 51172 1556 51224 1562
rect 51172 1498 51224 1504
rect 51184 800 51212 1498
rect 51264 1352 51316 1358
rect 51264 1294 51316 1300
rect 51276 898 51304 1294
rect 51350 1268 51410 2150
rect 55692 1970 55720 2751
rect 55784 2650 55812 3800
rect 55772 2644 55824 2650
rect 55772 2586 55824 2592
rect 55968 2582 55996 3800
rect 56230 3632 56286 3641
rect 56230 3567 56286 3576
rect 56046 3088 56102 3097
rect 56046 3023 56102 3032
rect 55956 2576 56008 2582
rect 55956 2518 56008 2524
rect 56060 2446 56088 3023
rect 56244 2650 56272 3567
rect 56336 3074 56364 3800
rect 56336 3046 56456 3074
rect 56428 2802 56456 3046
rect 56520 2990 56548 3800
rect 56600 3052 56652 3058
rect 56600 2994 56652 3000
rect 56508 2984 56560 2990
rect 56508 2926 56560 2932
rect 56612 2802 56640 2994
rect 56888 2922 56916 3800
rect 56876 2916 56928 2922
rect 56876 2858 56928 2864
rect 56428 2774 56640 2802
rect 57072 2650 57100 3800
rect 56232 2644 56284 2650
rect 56232 2586 56284 2592
rect 57060 2644 57112 2650
rect 57060 2586 57112 2592
rect 56324 2508 56376 2514
rect 56324 2450 56376 2456
rect 56048 2440 56100 2446
rect 56048 2382 56100 2388
rect 56230 2136 56286 2145
rect 56230 2071 56286 2080
rect 55864 2032 55916 2038
rect 55864 1974 55916 1980
rect 55954 2000 56010 2009
rect 55680 1964 55732 1970
rect 55680 1906 55732 1912
rect 55220 1896 55272 1902
rect 55220 1838 55272 1844
rect 53012 1556 53064 1562
rect 53012 1498 53064 1504
rect 51908 1488 51960 1494
rect 51908 1430 51960 1436
rect 52276 1488 52328 1494
rect 52276 1430 52328 1436
rect 52828 1488 52880 1494
rect 52828 1430 52880 1436
rect 51540 1420 51592 1426
rect 51592 1380 51764 1408
rect 51540 1362 51592 1368
rect 51350 1212 51352 1268
rect 51408 1212 51410 1268
rect 51350 1114 51410 1212
rect 51350 1062 51354 1114
rect 51406 1062 51410 1114
rect 51350 1040 51410 1062
rect 51276 870 51396 898
rect 51368 800 51396 870
rect 51736 800 51764 1380
rect 51920 800 51948 1430
rect 52288 800 52316 1430
rect 52460 1352 52512 1358
rect 52460 1294 52512 1300
rect 52472 800 52500 1294
rect 52840 800 52868 1430
rect 53024 800 53052 1498
rect 53656 1488 53708 1494
rect 54300 1488 54352 1494
rect 53708 1448 53788 1476
rect 53656 1430 53708 1436
rect 53288 1420 53340 1426
rect 53564 1420 53616 1426
rect 53340 1380 53420 1408
rect 53288 1362 53340 1368
rect 53392 800 53420 1380
rect 53564 1362 53616 1368
rect 53576 800 53604 1362
rect 53760 800 53788 1448
rect 54300 1430 54352 1436
rect 54852 1488 54904 1494
rect 54852 1430 54904 1436
rect 54116 1420 54168 1426
rect 54116 1362 54168 1368
rect 54128 800 54156 1362
rect 54312 800 54340 1430
rect 54668 1420 54720 1426
rect 54668 1362 54720 1368
rect 54680 800 54708 1362
rect 54864 800 54892 1430
rect 55232 800 55260 1838
rect 55588 1760 55640 1766
rect 55588 1702 55640 1708
rect 55404 1420 55456 1426
rect 55404 1362 55456 1368
rect 55416 800 55444 1362
rect 55600 800 55628 1702
rect 55876 1562 55904 1974
rect 56244 1970 56272 2071
rect 55954 1935 55956 1944
rect 56008 1935 56010 1944
rect 56232 1964 56284 1970
rect 55956 1906 56008 1912
rect 56232 1906 56284 1912
rect 55956 1828 56008 1834
rect 55956 1770 56008 1776
rect 55864 1556 55916 1562
rect 55864 1498 55916 1504
rect 55968 800 55996 1770
rect 56140 1284 56192 1290
rect 56140 1226 56192 1232
rect 56152 800 56180 1226
rect 56336 921 56364 2450
rect 57440 2446 57468 3800
rect 57624 2582 57652 3800
rect 57888 2916 57940 2922
rect 57992 2904 58020 3800
rect 58176 3058 58204 3800
rect 58360 3126 58388 3800
rect 58348 3120 58400 3126
rect 58348 3062 58400 3068
rect 58164 3052 58216 3058
rect 58164 2994 58216 3000
rect 57940 2876 58020 2904
rect 57888 2858 57940 2864
rect 57612 2576 57664 2582
rect 57612 2518 57664 2524
rect 57428 2440 57480 2446
rect 57428 2382 57480 2388
rect 58728 2378 58756 3800
rect 58912 3194 58940 3800
rect 58900 3188 58952 3194
rect 58900 3130 58952 3136
rect 59280 2854 59308 3800
rect 59268 2848 59320 2854
rect 59268 2790 59320 2796
rect 58716 2372 58768 2378
rect 58716 2314 58768 2320
rect 57980 2100 58032 2106
rect 57980 2042 58032 2048
rect 56784 1828 56836 1834
rect 56784 1770 56836 1776
rect 56508 1760 56560 1766
rect 56506 1728 56508 1737
rect 56600 1760 56652 1766
rect 56560 1728 56562 1737
rect 56600 1702 56652 1708
rect 56506 1663 56562 1672
rect 56508 1556 56560 1562
rect 56508 1498 56560 1504
rect 56322 912 56378 921
rect 56322 847 56378 856
rect 56520 800 56548 1498
rect 56612 1358 56640 1702
rect 56692 1420 56744 1426
rect 56692 1362 56744 1368
rect 56600 1352 56652 1358
rect 56600 1294 56652 1300
rect 56704 800 56732 1362
rect 56796 1057 56824 1770
rect 56980 1550 57284 1578
rect 56980 1494 57008 1550
rect 56968 1488 57020 1494
rect 56968 1430 57020 1436
rect 57060 1488 57112 1494
rect 57060 1430 57112 1436
rect 56782 1048 56838 1057
rect 56782 983 56838 992
rect 57072 800 57100 1430
rect 57256 800 57284 1550
rect 57612 1488 57664 1494
rect 57612 1430 57664 1436
rect 57624 800 57652 1430
rect 57796 1420 57848 1426
rect 57796 1362 57848 1368
rect 57808 800 57836 1362
rect 57992 800 58020 2042
rect 58532 2032 58584 2038
rect 58532 1974 58584 1980
rect 58348 1556 58400 1562
rect 58348 1498 58400 1504
rect 58360 800 58388 1498
rect 58544 800 58572 1974
rect 58900 1828 58952 1834
rect 58900 1770 58952 1776
rect 58912 800 58940 1770
rect 59084 1760 59136 1766
rect 59084 1702 59136 1708
rect 59096 800 59124 1702
rect 570 0 626 800
rect 754 0 810 800
rect 938 0 994 800
rect 1306 0 1362 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2594 0 2650 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 4986 0 5042 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9770 0 9826 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12162 0 12218 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14002 0 14058 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16394 0 16450 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18786 0 18842 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21178 0 21234 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23018 0 23074 800
rect 23386 0 23442 800
rect 23570 0 23626 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 24858 0 24914 800
rect 25226 0 25282 800
rect 25410 0 25466 800
rect 25778 0 25834 800
rect 25962 0 26018 800
rect 26146 0 26202 800
rect 26514 0 26570 800
rect 26698 0 26754 800
rect 27066 0 27122 800
rect 27250 0 27306 800
rect 27618 0 27674 800
rect 27802 0 27858 800
rect 27986 0 28042 800
rect 28354 0 28410 800
rect 28538 0 28594 800
rect 28906 0 28962 800
rect 29090 0 29146 800
rect 29458 0 29514 800
rect 29642 0 29698 800
rect 30010 0 30066 800
rect 30194 0 30250 800
rect 30378 0 30434 800
rect 30746 0 30802 800
rect 30930 0 30986 800
rect 31298 0 31354 800
rect 31482 0 31538 800
rect 31850 0 31906 800
rect 32034 0 32090 800
rect 32402 0 32458 800
rect 32586 0 32642 800
rect 32770 0 32826 800
rect 33138 0 33194 800
rect 33322 0 33378 800
rect 33690 0 33746 800
rect 33874 0 33930 800
rect 34242 0 34298 800
rect 34426 0 34482 800
rect 34794 0 34850 800
rect 34978 0 35034 800
rect 35162 0 35218 800
rect 35530 0 35586 800
rect 35714 0 35770 800
rect 36082 0 36138 800
rect 36266 0 36322 800
rect 36634 0 36690 800
rect 36818 0 36874 800
rect 37186 0 37242 800
rect 37370 0 37426 800
rect 37554 0 37610 800
rect 37922 0 37978 800
rect 38106 0 38162 800
rect 38474 0 38530 800
rect 38658 0 38714 800
rect 39026 0 39082 800
rect 39210 0 39266 800
rect 39578 0 39634 800
rect 39762 0 39818 800
rect 39946 0 40002 800
rect 40314 0 40370 800
rect 40498 0 40554 800
rect 40866 0 40922 800
rect 41050 0 41106 800
rect 41418 0 41474 800
rect 41602 0 41658 800
rect 41786 0 41842 800
rect 42154 0 42210 800
rect 42338 0 42394 800
rect 42706 0 42762 800
rect 42890 0 42946 800
rect 43258 0 43314 800
rect 43442 0 43498 800
rect 43810 0 43866 800
rect 43994 0 44050 800
rect 44178 0 44234 800
rect 44546 0 44602 800
rect 44730 0 44786 800
rect 45098 0 45154 800
rect 45282 0 45338 800
rect 45650 0 45706 800
rect 45834 0 45890 800
rect 46202 0 46258 800
rect 46386 0 46442 800
rect 46570 0 46626 800
rect 46938 0 46994 800
rect 47122 0 47178 800
rect 47490 0 47546 800
rect 47674 0 47730 800
rect 48042 0 48098 800
rect 48226 0 48282 800
rect 48594 0 48650 800
rect 48778 0 48834 800
rect 48962 0 49018 800
rect 49330 0 49386 800
rect 49514 0 49570 800
rect 49882 0 49938 800
rect 50066 0 50122 800
rect 50434 0 50490 800
rect 50618 0 50674 800
rect 50986 0 51042 800
rect 51170 0 51226 800
rect 51354 0 51410 800
rect 51722 0 51778 800
rect 51906 0 51962 800
rect 52274 0 52330 800
rect 52458 0 52514 800
rect 52826 0 52882 800
rect 53010 0 53066 800
rect 53378 0 53434 800
rect 53562 0 53618 800
rect 53746 0 53802 800
rect 54114 0 54170 800
rect 54298 0 54354 800
rect 54666 0 54722 800
rect 54850 0 54906 800
rect 55218 0 55274 800
rect 55402 0 55458 800
rect 55586 0 55642 800
rect 55954 0 56010 800
rect 56138 0 56194 800
rect 56506 0 56562 800
rect 56690 0 56746 800
rect 57058 0 57114 800
rect 57242 0 57298 800
rect 57610 0 57666 800
rect 57794 0 57850 800
rect 57978 0 58034 800
rect 58346 0 58402 800
rect 58530 0 58586 800
rect 58898 0 58954 800
rect 59082 0 59138 800
<< via2 >>
rect 3146 3576 3202 3632
rect 3974 3032 4030 3088
rect 4158 2760 4214 2816
rect 2870 992 2926 1048
rect 3974 2080 4030 2136
rect 3698 1964 3754 2000
rect 3698 1944 3700 1964
rect 3700 1944 3752 1964
rect 3752 1944 3754 1964
rect 11352 2292 11408 2348
rect 3514 1420 3570 1456
rect 3514 1400 3516 1420
rect 3516 1400 3568 1420
rect 3568 1400 3570 1420
rect 3352 1212 3408 1268
rect 19352 1212 19408 1268
rect 25502 2488 25558 2544
rect 23294 1980 23296 2000
rect 23296 1980 23348 2000
rect 23348 1980 23350 2000
rect 23294 1944 23350 1980
rect 25226 1944 25282 2000
rect 25042 1556 25098 1592
rect 25042 1536 25044 1556
rect 25044 1536 25096 1556
rect 25096 1536 25098 1556
rect 26146 2524 26148 2544
rect 26148 2524 26200 2544
rect 26200 2524 26202 2544
rect 25962 1536 26018 1592
rect 26146 2488 26202 2524
rect 27352 2292 27408 2348
rect 43352 2292 43408 2348
rect 35352 1212 35408 1268
rect 55678 2760 55734 2816
rect 56230 3576 56286 3632
rect 56046 3032 56102 3088
rect 56230 2080 56286 2136
rect 51352 1212 51408 1268
rect 55954 1964 56010 2000
rect 55954 1944 55956 1964
rect 55956 1944 56008 1964
rect 56008 1944 56010 1964
rect 56506 1708 56508 1728
rect 56508 1708 56560 1728
rect 56560 1708 56562 1728
rect 56506 1672 56562 1708
rect 56322 856 56378 912
rect 56782 992 56838 1048
<< metal3 >>
rect 0 3634 800 3664
rect 3141 3634 3207 3637
rect 0 3632 3207 3634
rect 0 3576 3146 3632
rect 3202 3576 3207 3632
rect 0 3574 3207 3576
rect 0 3544 800 3574
rect 3141 3571 3207 3574
rect 56225 3634 56291 3637
rect 59200 3634 60000 3664
rect 56225 3632 60000 3634
rect 56225 3576 56230 3632
rect 56286 3576 60000 3632
rect 56225 3574 60000 3576
rect 56225 3571 56291 3574
rect 59200 3544 60000 3574
rect 0 3090 800 3120
rect 3969 3090 4035 3093
rect 0 3088 4035 3090
rect 0 3032 3974 3088
rect 4030 3032 4035 3088
rect 0 3030 4035 3032
rect 0 3000 800 3030
rect 3969 3027 4035 3030
rect 56041 3090 56107 3093
rect 59200 3090 60000 3120
rect 56041 3088 60000 3090
rect 56041 3032 56046 3088
rect 56102 3032 60000 3088
rect 56041 3030 60000 3032
rect 56041 3027 56107 3030
rect 59200 3000 60000 3030
rect 0 2818 800 2848
rect 4153 2818 4219 2821
rect 0 2816 4219 2818
rect 0 2760 4158 2816
rect 4214 2760 4219 2816
rect 0 2758 4219 2760
rect 0 2728 800 2758
rect 4153 2755 4219 2758
rect 55673 2818 55739 2821
rect 59200 2818 60000 2848
rect 55673 2816 60000 2818
rect 55673 2760 55678 2816
rect 55734 2760 60000 2816
rect 55673 2758 60000 2760
rect 55673 2755 55739 2758
rect 59200 2728 60000 2758
rect 25497 2546 25563 2549
rect 26141 2546 26207 2549
rect 25497 2544 26207 2546
rect 25497 2488 25502 2544
rect 25558 2488 26146 2544
rect 26202 2488 26207 2544
rect 25497 2486 26207 2488
rect 25497 2483 25563 2486
rect 26141 2483 26207 2486
rect 11347 2350 11413 2353
rect 27347 2350 27413 2353
rect 43347 2350 43413 2353
rect 1380 2348 58604 2350
rect 0 2274 800 2304
rect 1380 2292 11352 2348
rect 11408 2292 27352 2348
rect 27408 2292 43352 2348
rect 43408 2292 58604 2348
rect 1380 2290 58604 2292
rect 11347 2287 11413 2290
rect 27347 2287 27413 2290
rect 43347 2287 43413 2290
rect 59200 2274 60000 2304
rect 0 2214 1226 2274
rect 0 2184 800 2214
rect 1166 2138 1226 2214
rect 58758 2214 60000 2274
rect 3969 2138 4035 2141
rect 1166 2136 4035 2138
rect 1166 2080 3974 2136
rect 4030 2080 4035 2136
rect 1166 2078 4035 2080
rect 3969 2075 4035 2078
rect 56225 2138 56291 2141
rect 58758 2138 58818 2214
rect 59200 2184 60000 2214
rect 56225 2136 58818 2138
rect 56225 2080 56230 2136
rect 56286 2080 58818 2136
rect 56225 2078 58818 2080
rect 56225 2075 56291 2078
rect 0 2002 800 2032
rect 3693 2002 3759 2005
rect 0 2000 3759 2002
rect 0 1944 3698 2000
rect 3754 1944 3759 2000
rect 0 1942 3759 1944
rect 0 1912 800 1942
rect 3693 1939 3759 1942
rect 23289 2002 23355 2005
rect 25221 2002 25287 2005
rect 23289 2000 25287 2002
rect 23289 1944 23294 2000
rect 23350 1944 25226 2000
rect 25282 1944 25287 2000
rect 23289 1942 25287 1944
rect 23289 1939 23355 1942
rect 25221 1939 25287 1942
rect 55949 2002 56015 2005
rect 59200 2002 60000 2032
rect 55949 2000 60000 2002
rect 55949 1944 55954 2000
rect 56010 1944 60000 2000
rect 55949 1942 60000 1944
rect 55949 1939 56015 1942
rect 59200 1912 60000 1942
rect 56501 1730 56567 1733
rect 59200 1730 60000 1760
rect 56501 1728 60000 1730
rect 56501 1672 56506 1728
rect 56562 1672 60000 1728
rect 56501 1670 60000 1672
rect 56501 1667 56567 1670
rect 59200 1640 60000 1670
rect 25037 1594 25103 1597
rect 25957 1594 26023 1597
rect 25037 1592 26023 1594
rect 25037 1536 25042 1592
rect 25098 1536 25962 1592
rect 26018 1536 26023 1592
rect 25037 1534 26023 1536
rect 25037 1531 25103 1534
rect 25957 1531 26023 1534
rect 0 1458 800 1488
rect 3509 1458 3575 1461
rect 0 1456 3575 1458
rect 0 1400 3514 1456
rect 3570 1400 3575 1456
rect 0 1398 3575 1400
rect 0 1368 800 1398
rect 3509 1395 3575 1398
rect 3347 1270 3413 1273
rect 19347 1270 19413 1273
rect 35347 1270 35413 1273
rect 51347 1270 51413 1273
rect 1380 1268 58604 1270
rect 0 1186 800 1216
rect 1380 1212 3352 1268
rect 3408 1212 19352 1268
rect 19408 1212 35352 1268
rect 35408 1212 51352 1268
rect 51408 1212 58604 1268
rect 1380 1210 58604 1212
rect 3347 1207 3413 1210
rect 19347 1207 19413 1210
rect 35347 1207 35413 1210
rect 51347 1207 51413 1210
rect 59200 1186 60000 1216
rect 0 1126 1226 1186
rect 0 1096 800 1126
rect 1166 1050 1226 1126
rect 58758 1126 60000 1186
rect 2865 1050 2931 1053
rect 1166 1048 2931 1050
rect 1166 992 2870 1048
rect 2926 992 2931 1048
rect 1166 990 2931 992
rect 2865 987 2931 990
rect 56777 1050 56843 1053
rect 58758 1050 58818 1126
rect 59200 1096 60000 1126
rect 56777 1048 58818 1050
rect 56777 992 56782 1048
rect 56838 992 58818 1048
rect 56777 990 58818 992
rect 56777 987 56843 990
rect 56317 914 56383 917
rect 59200 914 60000 944
rect 56317 912 60000 914
rect 56317 856 56322 912
rect 56378 856 60000 912
rect 56317 854 60000 856
rect 56317 851 56383 854
rect 59200 824 60000 854
use sky130_fd_sc_hd__conb_1  insts\[42\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607116009
transform 1 0 2300 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[449\]
timestamp 1607116009
transform 1 0 2024 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607116009
transform 1 0 1380 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1607116009
transform 1 0 1380 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607116009
transform 1 0 1656 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607116009
transform 1 0 1656 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607116009
transform 1 0 2760 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[411\]
timestamp 1607116009
transform 1 0 2576 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[371\]
timestamp 1607116009
transform 1 0 2852 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[268\]
timestamp 1607116009
transform 1 0 2852 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[321\]
timestamp 1607116009
transform 1 0 3128 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[221\]
timestamp 1607116009
transform 1 0 3128 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[301\]
timestamp 1607116009
transform 1 0 3404 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[213\]
timestamp 1607116009
transform 1 0 3404 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[201\]
timestamp 1607116009
transform 1 0 3680 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[105\]
timestamp 1607116009
transform 1 0 3680 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[110\]
timestamp 1607116009
transform 1 0 3956 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[176\]
timestamp 1607116009
transform 1 0 4324 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[223\]
timestamp 1607116009
transform 1 0 3956 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[235\]
timestamp 1607116009
transform 1 0 4600 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[240\]
timestamp 1607116009
transform 1 0 4876 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[258\]
timestamp 1607116009
transform 1 0 4508 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[270\]
timestamp 1607116009
transform 1 0 4232 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[43\]
timestamp 1607116009
transform 1 0 4784 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607116009
transform 1 0 4232 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[116\]
timestamp 1607116009
transform 1 0 5980 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[177\]
timestamp 1607116009
transform 1 0 5336 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[346\]
timestamp 1607116009
transform 1 0 5612 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[388\]
timestamp 1607116009
transform 1 0 5612 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[68\]
timestamp 1607116009
transform 1 0 5060 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[71\]
timestamp 1607116009
transform 1 0 5336 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607116009
transform 1 0 5152 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49
timestamp 1607116009
transform 1 0 5888 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_49
timestamp 1607116009
transform 1 0 5888 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[180\]
timestamp 1607116009
transform 1 0 6256 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[26\]
timestamp 1607116009
transform 1 0 6624 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[320\]
timestamp 1607116009
transform 1 0 7176 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_9
timestamp 1607116009
transform 1 0 7084 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_27
timestamp 1607116009
transform 1 0 6992 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56
timestamp 1607116009
transform 1 0 6532 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1607116009
transform 1 0 6900 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_62 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607116009
transform 1 0 7084 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[12\]
timestamp 1607116009
transform 1 0 8188 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[143\]
timestamp 1607116009
transform 1 0 7544 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[159\]
timestamp 1607116009
transform 1 0 8464 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[323\]
timestamp 1607116009
transform 1 0 7820 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[47\]
timestamp 1607116009
transform 1 0 8004 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66
timestamp 1607116009
transform 1 0 7452 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73
timestamp 1607116009
transform 1 0 8096 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_70
timestamp 1607116009
transform 1 0 7820 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_75
timestamp 1607116009
transform 1 0 8280 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[219\]
timestamp 1607116009
transform 1 0 8740 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[310\]
timestamp 1607116009
transform 1 0 9016 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[317\]
timestamp 1607116009
transform 1 0 9568 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[362\]
timestamp 1607116009
transform 1 0 9292 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_87
timestamp 1607116009
transform 1 0 9384 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[112\]
timestamp 1607116009
transform 1 0 10212 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[139\]
timestamp 1607116009
transform 1 0 10488 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[185\]
timestamp 1607116009
transform 1 0 10580 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_10
timestamp 1607116009
transform 1 0 9936 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 1607116009
transform 1 0 9844 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_94
timestamp 1607116009
transform 1 0 10028 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_102
timestamp 1607116009
transform 1 0 10764 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_99
timestamp 1607116009
transform 1 0 10488 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_107
timestamp 1607116009
transform 1 0 11224 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_103
timestamp 1607116009
transform 1 0 10856 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  insts\[168\]
timestamp 1607116009
transform 1 0 11224 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[106\]
timestamp 1607116009
transform 1 0 10948 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_111
timestamp 1607116009
transform 1 0 11592 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  insts\[448\]
timestamp 1607116009
transform 1 0 11316 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[187\]
timestamp 1607116009
transform 1 0 11500 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_115
timestamp 1607116009
transform 1 0 11960 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113
timestamp 1607116009
transform 1 0 11776 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[119\]
timestamp 1607116009
transform 1 0 11868 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_119
timestamp 1607116009
transform 1 0 12328 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117
timestamp 1607116009
transform 1 0 12144 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[314\]
timestamp 1607116009
transform 1 0 12052 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[149\]
timestamp 1607116009
transform 1 0 12328 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1607116009
transform 1 0 12604 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_28
timestamp 1607116009
transform 1 0 12604 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[181\]
timestamp 1607116009
transform 1 0 12696 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_11
timestamp 1607116009
transform 1 0 12788 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[231\]
timestamp 1607116009
transform 1 0 12972 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[115\]
timestamp 1607116009
transform 1 0 12880 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[170\]
timestamp 1607116009
transform 1 0 13156 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[160\]
timestamp 1607116009
transform 1 0 13984 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[1\]
timestamp 1607116009
transform 1 0 13432 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[232\]
timestamp 1607116009
transform 1 0 13708 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[331\]
timestamp 1607116009
transform 1 0 14260 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[397\]
timestamp 1607116009
transform 1 0 13248 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[413\]
timestamp 1607116009
transform 1 0 13524 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[62\]
timestamp 1607116009
transform 1 0 13800 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_138
timestamp 1607116009
transform 1 0 14076 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  insts\[249\]
timestamp 1607116009
transform 1 0 14628 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[265\]
timestamp 1607116009
transform 1 0 14996 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[324\]
timestamp 1607116009
transform 1 0 15272 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[379\]
timestamp 1607116009
transform 1 0 14444 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_143
timestamp 1607116009
transform 1 0 14536 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_147
timestamp 1607116009
transform 1 0 14904 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1607116009
transform 1 0 15548 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_145
timestamp 1607116009
transform 1 0 14720 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[251\]
timestamp 1607116009
transform 1 0 16652 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[341\]
timestamp 1607116009
transform 1 0 15732 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[378\]
timestamp 1607116009
transform 1 0 16008 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[3\]
timestamp 1607116009
transform 1 0 16376 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_12
timestamp 1607116009
transform 1 0 15640 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_162
timestamp 1607116009
transform 1 0 16284 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_157
timestamp 1607116009
transform 1 0 15824 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[212\]
timestamp 1607116009
transform 1 0 17756 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[245\]
timestamp 1607116009
transform 1 0 17296 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[414\]
timestamp 1607116009
transform 1 0 16928 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[436\]
timestamp 1607116009
transform 1 0 17020 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_172
timestamp 1607116009
transform 1 0 17204 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_176
timestamp 1607116009
transform 1 0 17572 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_169
timestamp 1607116009
transform 1 0 16928 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_173
timestamp 1607116009
transform 1 0 17296 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_184
timestamp 1607116009
transform 1 0 18308 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1607116009
transform 1 0 18032 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1607116009
transform 1 0 18308 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_29
timestamp 1607116009
transform 1 0 18216 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_13
timestamp 1607116009
transform 1 0 18492 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[96\]
timestamp 1607116009
transform 1 0 18032 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_190
timestamp 1607116009
transform 1 0 18860 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[437\]
timestamp 1607116009
transform 1 0 18584 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[293\]
timestamp 1607116009
transform 1 0 19044 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[129\]
timestamp 1607116009
transform 1 0 18584 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_190
timestamp 1607116009
transform 1 0 18860 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[211\]
timestamp 1607116009
transform 1 0 20056 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[311\]
timestamp 1607116009
transform 1 0 19412 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[349\]
timestamp 1607116009
transform 1 0 19688 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1607116009
transform 1 0 19320 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_202
timestamp 1607116009
transform 1 0 19964 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_202
timestamp 1607116009
transform 1 0 19964 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[386\]
timestamp 1607116009
transform 1 0 20608 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[373\]
timestamp 1607116009
transform 1 0 20332 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_210
timestamp 1607116009
transform 1 0 20700 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[66\]
timestamp 1607116009
transform 1 0 20792 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[40\]
timestamp 1607116009
transform 1 0 20884 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1607116009
transform 1 0 21160 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[64\]
timestamp 1607116009
transform 1 0 21068 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_14
timestamp 1607116009
transform 1 0 21344 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[289\]
timestamp 1607116009
transform 1 0 21344 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[22\]
timestamp 1607116009
transform 1 0 21436 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[103\]
timestamp 1607116009
transform 1 0 22264 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[15\]
timestamp 1607116009
transform 1 0 22540 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[399\]
timestamp 1607116009
transform 1 0 22172 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[440\]
timestamp 1607116009
transform 1 0 21896 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[447\]
timestamp 1607116009
transform 1 0 22448 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[56\]
timestamp 1607116009
transform 1 0 21896 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[61\]
timestamp 1607116009
transform 1 0 21620 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1607116009
transform 1 0 21712 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_226
timestamp 1607116009
transform 1 0 22172 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1607116009
transform 1 0 22816 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[391\]
timestamp 1607116009
transform 1 0 22724 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[156\]
timestamp 1607116009
transform 1 0 22908 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_235
timestamp 1607116009
transform 1 0 23000 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_237
timestamp 1607116009
transform 1 0 23184 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[392\]
timestamp 1607116009
transform 1 0 23092 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_242
timestamp 1607116009
transform 1 0 23644 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_242
timestamp 1607116009
transform 1 0 23644 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[200\]
timestamp 1607116009
transform 1 0 23368 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[125\]
timestamp 1607116009
transform 1 0 23368 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[17\]
timestamp 1607116009
transform 1 0 23736 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_245
timestamp 1607116009
transform 1 0 23920 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_246
timestamp 1607116009
transform 1 0 24012 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_30
timestamp 1607116009
transform 1 0 23828 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[254\]
timestamp 1607116009
transform 1 0 24012 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_15
timestamp 1607116009
transform 1 0 24196 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[318\]
timestamp 1607116009
transform 1 0 24288 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[166\]
timestamp 1607116009
transform 1 0 24288 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_252
timestamp 1607116009
transform 1 0 24564 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[344\]
timestamp 1607116009
transform 1 0 24748 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[214\]
timestamp 1607116009
transform 1 0 24840 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[202\]
timestamp 1607116009
transform 1 0 24564 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[452\]
timestamp 1607116009
transform 1 0 25024 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[330\]
timestamp 1607116009
transform 1 0 25300 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[302\]
timestamp 1607116009
transform 1 0 25116 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_264
timestamp 1607116009
transform 1 0 25668 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[365\]
timestamp 1607116009
transform 1 0 25576 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[327\]
timestamp 1607116009
transform 1 0 25392 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[36\]
timestamp 1607116009
transform 1 0 25852 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[329\]
timestamp 1607116009
transform 1 0 26036 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[150\]
timestamp 1607116009
transform 1 0 25760 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[382\]
timestamp 1607116009
transform 1 0 26128 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[157\]
timestamp 1607116009
transform 1 0 27140 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[199\]
timestamp 1607116009
transform 1 0 26312 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[415\]
timestamp 1607116009
transform 1 0 26588 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[93\]
timestamp 1607116009
transform 1 0 26404 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_16
timestamp 1607116009
transform 1 0 27048 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_277
timestamp 1607116009
transform 1 0 26864 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_275
timestamp 1607116009
transform 1 0 26680 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[220\]
timestamp 1607116009
transform 1 0 27692 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[23\]
timestamp 1607116009
transform 1 0 28336 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[284\]
timestamp 1607116009
transform 1 0 27416 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[419\]
timestamp 1607116009
transform 1 0 27968 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[455\]
timestamp 1607116009
transform 1 0 27968 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_292
timestamp 1607116009
transform 1 0 28244 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_287
timestamp 1607116009
transform 1 0 27784 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_292
timestamp 1607116009
transform 1 0 28244 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[326\]
timestamp 1607116009
transform 1 0 29164 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[39\]
timestamp 1607116009
transform 1 0 28612 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[400\]
timestamp 1607116009
transform 1 0 29532 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[446\]
timestamp 1607116009
transform 1 0 28888 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_31
timestamp 1607116009
transform 1 0 29440 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_305
timestamp 1607116009
transform 1 0 29440 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_304
timestamp 1607116009
transform 1 0 29348 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_306
timestamp 1607116009
transform 1 0 29532 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[171\]
timestamp 1607116009
transform 1 0 30636 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[315\]
timestamp 1607116009
transform 1 0 29992 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[334\]
timestamp 1607116009
transform 1 0 30268 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[67\]
timestamp 1607116009
transform 1 0 30360 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_17
timestamp 1607116009
transform 1 0 29900 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_309
timestamp 1607116009
transform 1 0 29808 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_317
timestamp 1607116009
transform 1 0 30544 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_314
timestamp 1607116009
transform 1 0 30268 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_318
timestamp 1607116009
transform 1 0 30636 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  insts\[132\]
timestamp 1607116009
transform 1 0 31188 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[278\]
timestamp 1607116009
transform 1 0 31556 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[351\]
timestamp 1607116009
transform 1 0 31832 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[420\]
timestamp 1607116009
transform 1 0 30912 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[86\]
timestamp 1607116009
transform 1 0 31096 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_327
timestamp 1607116009
transform 1 0 31464 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_322
timestamp 1607116009
transform 1 0 31004 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_326
timestamp 1607116009
transform 1 0 31372 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[102\]
timestamp 1607116009
transform 1 0 33212 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[142\]
timestamp 1607116009
transform 1 0 32200 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[172\]
timestamp 1607116009
transform 1 0 32476 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[424\]
timestamp 1607116009
transform 1 0 32844 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_18
timestamp 1607116009
transform 1 0 32752 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_334
timestamp 1607116009
transform 1 0 32108 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_345
timestamp 1607116009
transform 1 0 33120 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_338
timestamp 1607116009
transform 1 0 32476 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[14\]
timestamp 1607116009
transform 1 0 33580 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[283\]
timestamp 1607116009
transform 1 0 34408 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[401\]
timestamp 1607116009
transform 1 0 34132 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[417\]
timestamp 1607116009
transform 1 0 33856 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[9\]
timestamp 1607116009
transform 1 0 33856 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_349
timestamp 1607116009
transform 1 0 33488 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_350
timestamp 1607116009
transform 1 0 33580 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_356
timestamp 1607116009
transform 1 0 34132 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[208\]
timestamp 1607116009
transform 1 0 35052 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[299\]
timestamp 1607116009
transform 1 0 35328 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[305\]
timestamp 1607116009
transform 1 0 34776 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_19
timestamp 1607116009
transform 1 0 35604 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_32
timestamp 1607116009
transform 1 0 35052 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_362
timestamp 1607116009
transform 1 0 34684 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_364
timestamp 1607116009
transform 1 0 34868 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_367
timestamp 1607116009
transform 1 0 35144 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[182\]
timestamp 1607116009
transform 1 0 36800 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[195\]
timestamp 1607116009
transform 1 0 36432 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[266\]
timestamp 1607116009
transform 1 0 35696 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[28\]
timestamp 1607116009
transform 1 0 35972 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_379
timestamp 1607116009
transform 1 0 36248 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_384
timestamp 1607116009
transform 1 0 36708 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_379
timestamp 1607116009
transform 1 0 36248 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[215\]
timestamp 1607116009
transform 1 0 37628 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[303\]
timestamp 1607116009
transform 1 0 37904 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[345\]
timestamp 1607116009
transform 1 0 37904 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[410\]
timestamp 1607116009
transform 1 0 37076 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[4\]
timestamp 1607116009
transform 1 0 37352 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_391 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607116009
transform 1 0 37352 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  insts\[222\]
timestamp 1607116009
transform 1 0 38548 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[276\]
timestamp 1607116009
transform 1 0 38916 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[296\]
timestamp 1607116009
transform 1 0 38180 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_20
timestamp 1607116009
transform 1 0 38456 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_407
timestamp 1607116009
transform 1 0 38824 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_400
timestamp 1607116009
transform 1 0 38180 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[120\]
timestamp 1607116009
transform 1 0 39836 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[297\]
timestamp 1607116009
transform 1 0 40204 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[30\]
timestamp 1607116009
transform 1 0 39560 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[405\]
timestamp 1607116009
transform 1 0 39192 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[69\]
timestamp 1607116009
transform 1 0 39468 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_414
timestamp 1607116009
transform 1 0 39468 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_421
timestamp 1607116009
transform 1 0 40112 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_412
timestamp 1607116009
transform 1 0 39284 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_417
timestamp 1607116009
transform 1 0 39744 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_428
timestamp 1607116009
transform 1 0 40756 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_425
timestamp 1607116009
transform 1 0 40480 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_428
timestamp 1607116009
transform 1 0 40756 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_33
timestamp 1607116009
transform 1 0 40664 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[216\]
timestamp 1607116009
transform 1 0 40480 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[108\]
timestamp 1607116009
transform 1 0 40848 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_435
timestamp 1607116009
transform 1 0 41400 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_432
timestamp 1607116009
transform 1 0 41124 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_21
timestamp 1607116009
transform 1 0 41308 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[319\]
timestamp 1607116009
transform 1 0 41124 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[153\]
timestamp 1607116009
transform 1 0 41492 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_435
timestamp 1607116009
transform 1 0 41400 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[237\]
timestamp 1607116009
transform 1 0 41768 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[34\]
timestamp 1607116009
transform 1 0 42136 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[394\]
timestamp 1607116009
transform 1 0 42504 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[407\]
timestamp 1607116009
transform 1 0 42320 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_442
timestamp 1607116009
transform 1 0 42044 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_446
timestamp 1607116009
transform 1 0 42412 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_443
timestamp 1607116009
transform 1 0 42136 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_448
timestamp 1607116009
transform 1 0 42596 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  insts\[209\]
timestamp 1607116009
transform 1 0 43700 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[277\]
timestamp 1607116009
transform 1 0 43424 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[307\]
timestamp 1607116009
transform 1 0 42964 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[428\]
timestamp 1607116009
transform 1 0 43148 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_450
timestamp 1607116009
transform 1 0 42780 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_455
timestamp 1607116009
transform 1 0 43240 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_457
timestamp 1607116009
transform 1 0 43424 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[114\]
timestamp 1607116009
transform 1 0 44896 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[228\]
timestamp 1607116009
transform 1 0 44344 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[458\]
timestamp 1607116009
transform 1 0 44620 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_22
timestamp 1607116009
transform 1 0 44160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_463
timestamp 1607116009
transform 1 0 43976 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_466
timestamp 1607116009
transform 1 0 44252 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_469
timestamp 1607116009
transform 1 0 44528 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  insts\[175\]
timestamp 1607116009
transform 1 0 46184 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[204\]
timestamp 1607116009
transform 1 0 45724 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[29\]
timestamp 1607116009
transform 1 0 45172 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[367\]
timestamp 1607116009
transform 1 0 45448 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[6\]
timestamp 1607116009
transform 1 0 45172 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_485
timestamp 1607116009
transform 1 0 46000 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_475
timestamp 1607116009
transform 1 0 45080 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_479
timestamp 1607116009
transform 1 0 45448 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_487
timestamp 1607116009
transform 1 0 46184 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[280\]
timestamp 1607116009
transform 1 0 47104 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[31\]
timestamp 1607116009
transform 1 0 46460 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[63\]
timestamp 1607116009
transform 1 0 46736 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_23
timestamp 1607116009
transform 1 0 47012 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_34
timestamp 1607116009
transform 1 0 46276 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_500
timestamp 1607116009
transform 1 0 47380 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_489
timestamp 1607116009
transform 1 0 46368 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[255\]
timestamp 1607116009
transform 1 0 47472 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[360\]
timestamp 1607116009
transform 1 0 48116 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[406\]
timestamp 1607116009
transform 1 0 47748 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[456\]
timestamp 1607116009
transform 1 0 48392 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[7\]
timestamp 1607116009
transform 1 0 48300 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_507
timestamp 1607116009
transform 1 0 48024 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_501
timestamp 1607116009
transform 1 0 47472 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_509
timestamp 1607116009
transform 1 0 48208 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_513
timestamp 1607116009
transform 1 0 48576 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[13\]
timestamp 1607116009
transform 1 0 49312 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[234\]
timestamp 1607116009
transform 1 0 48668 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[295\]
timestamp 1607116009
transform 1 0 48944 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[384\]
timestamp 1607116009
transform 1 0 49588 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_520
timestamp 1607116009
transform 1 0 49220 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_525
timestamp 1607116009
transform 1 0 49680 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[261\]
timestamp 1607116009
transform 1 0 50140 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[369\]
timestamp 1607116009
transform 1 0 50416 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[46\]
timestamp 1607116009
transform 1 0 50784 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[65\]
timestamp 1607116009
transform 1 0 49956 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_24
timestamp 1607116009
transform 1 0 49864 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_528
timestamp 1607116009
transform 1 0 49956 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_536
timestamp 1607116009
transform 1 0 50692 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_531
timestamp 1607116009
transform 1 0 50232 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[203\]
timestamp 1607116009
transform 1 0 51336 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[264\]
timestamp 1607116009
transform 1 0 51612 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[48\]
timestamp 1607116009
transform 1 0 51060 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_35
timestamp 1607116009
transform 1 0 51888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_549
timestamp 1607116009
transform 1 0 51888 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_543
timestamp 1607116009
transform 1 0 51336 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_550
timestamp 1607116009
transform 1 0 51980 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[190\]
timestamp 1607116009
transform 1 0 52164 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[262\]
timestamp 1607116009
transform 1 0 52808 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[313\]
timestamp 1607116009
transform 1 0 53084 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[59\]
timestamp 1607116009
transform 1 0 52440 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_25
timestamp 1607116009
transform 1 0 52716 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_562
timestamp 1607116009
transform 1 0 53084 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[10\]
timestamp 1607116009
transform 1 0 54372 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[239\]
timestamp 1607116009
transform 1 0 53728 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[246\]
timestamp 1607116009
transform 1 0 54004 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[343\]
timestamp 1607116009
transform 1 0 53360 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[82\]
timestamp 1607116009
transform 1 0 54464 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_568
timestamp 1607116009
transform 1 0 53636 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_575
timestamp 1607116009
transform 1 0 54280 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_574
timestamp 1607116009
transform 1 0 54188 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[368\]
timestamp 1607116009
transform 1 0 54740 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[194\]
timestamp 1607116009
transform 1 0 54648 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_583
timestamp 1607116009
transform 1 0 55016 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_585
timestamp 1607116009
transform 1 0 55200 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[412\]
timestamp 1607116009
transform 1 0 55200 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[279\]
timestamp 1607116009
transform 1 0 54924 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_588
timestamp 1607116009
transform 1 0 55476 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_26
timestamp 1607116009
transform 1 0 55568 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[357\]
timestamp 1607116009
transform 1 0 55292 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[439\]
timestamp 1607116009
transform 1 0 55660 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[335\]
timestamp 1607116009
transform 1 0 55660 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[100\]
timestamp 1607116009
transform 1 0 55936 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[158\]
timestamp 1607116009
transform 1 0 55936 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[198\]
timestamp 1607116009
transform 1 0 56212 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[20\]
timestamp 1607116009
transform 1 0 56488 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[285\]
timestamp 1607116009
transform 1 0 56212 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[294\]
timestamp 1607116009
transform 1 0 56764 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[361\]
timestamp 1607116009
transform 1 0 56488 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[363\]
timestamp 1607116009
transform 1 0 56764 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[390\]
timestamp 1607116009
transform 1 0 57040 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[423\]
timestamp 1607116009
transform 1 0 57316 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[451\]
timestamp 1607116009
transform 1 0 57040 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[50\]
timestamp 1607116009
transform 1 0 57592 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[51\]
timestamp 1607116009
transform 1 0 57868 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[55\]
timestamp 1607116009
transform 1 0 57592 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_36
timestamp 1607116009
transform 1 0 57500 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_608
timestamp 1607116009
transform 1 0 57316 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_614
timestamp 1607116009
transform 1 0 57868 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1607116009
transform -1 0 58604 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1607116009
transform -1 0 58604 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_617
timestamp 1607116009
transform 1 0 58144 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_618
timestamp 1607116009
transform 1 0 58236 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1607116009
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1607116009
transform 1 0 1656 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[225\]
timestamp 1607116009
transform 1 0 3680 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[381\]
timestamp 1607116009
transform 1 0 3404 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[429\]
timestamp 1607116009
transform 1 0 3128 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[89\]
timestamp 1607116009
transform 1 0 2852 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_15
timestamp 1607116009
transform 1 0 2760 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[281\]
timestamp 1607116009
transform 1 0 3956 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[33\]
timestamp 1607116009
transform 1 0 4324 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[72\]
timestamp 1607116009
transform 1 0 4600 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[92\]
timestamp 1607116009
transform 1 0 4876 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_37
timestamp 1607116009
transform 1 0 4232 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1607116009
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1607116009
transform 1 0 6256 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1607116009
transform 1 0 7360 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1607116009
transform 1 0 8464 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  insts\[44\]
timestamp 1607116009
transform 1 0 9108 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1607116009
transform 1 0 9016 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_87
timestamp 1607116009
transform 1 0 9384 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_38
timestamp 1607116009
transform 1 0 9844 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1607116009
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1607116009
transform 1 0 9936 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[85\]
timestamp 1607116009
transform 1 0 11132 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_105
timestamp 1607116009
transform 1 0 11040 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_109
timestamp 1607116009
transform 1 0 11408 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[422\]
timestamp 1607116009
transform 1 0 13064 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_121
timestamp 1607116009
transform 1 0 12512 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_130
timestamp 1607116009
transform 1 0 13340 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_39
timestamp 1607116009
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_142
timestamp 1607116009
transform 1 0 14444 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_150
timestamp 1607116009
transform 1 0 15180 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1607116009
transform 1 0 15548 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_166
timestamp 1607116009
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[97\]
timestamp 1607116009
transform 1 0 16836 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_171
timestamp 1607116009
transform 1 0 17112 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[83\]
timestamp 1607116009
transform 1 0 18952 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_183
timestamp 1607116009
transform 1 0 18216 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[457\]
timestamp 1607116009
transform 1 0 19320 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_194
timestamp 1607116009
transform 1 0 19228 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_198
timestamp 1607116009
transform 1 0 19596 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[178\]
timestamp 1607116009
transform 1 0 20792 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[25\]
timestamp 1607116009
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[372\]
timestamp 1607116009
transform 1 0 20516 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_40
timestamp 1607116009
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_206
timestamp 1607116009
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_218
timestamp 1607116009
transform 1 0 21436 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[191\]
timestamp 1607116009
transform 1 0 21988 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[263\]
timestamp 1607116009
transform 1 0 21528 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[38\]
timestamp 1607116009
transform 1 0 22448 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_222
timestamp 1607116009
transform 1 0 21804 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_227
timestamp 1607116009
transform 1 0 22264 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[197\]
timestamp 1607116009
transform 1 0 22724 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[207\]
timestamp 1607116009
transform 1 0 23552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[325\]
timestamp 1607116009
transform 1 0 23184 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_235
timestamp 1607116009
transform 1 0 23000 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_240
timestamp 1607116009
transform 1 0 23460 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[184\]
timestamp 1607116009
transform 1 0 24288 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[287\]
timestamp 1607116009
transform 1 0 24932 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[342\]
timestamp 1607116009
transform 1 0 24656 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[348\]
timestamp 1607116009
transform 1 0 23828 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_247
timestamp 1607116009
transform 1 0 24104 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_252
timestamp 1607116009
transform 1 0 24564 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[253\]
timestamp 1607116009
transform 1 0 25392 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[267\]
timestamp 1607116009
transform 1 0 25852 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_259
timestamp 1607116009
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_264
timestamp 1607116009
transform 1 0 25668 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_269
timestamp 1607116009
transform 1 0 26128 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[146\]
timestamp 1607116009
transform 1 0 26220 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[282\]
timestamp 1607116009
transform 1 0 27048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[375\]
timestamp 1607116009
transform 1 0 26772 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[91\]
timestamp 1607116009
transform 1 0 27324 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_41
timestamp 1607116009
transform 1 0 26680 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_273
timestamp 1607116009
transform 1 0 26496 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[101\]
timestamp 1607116009
transform 1 0 28336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[21\]
timestamp 1607116009
transform 1 0 27692 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[272\]
timestamp 1607116009
transform 1 0 27968 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_285
timestamp 1607116009
transform 1 0 27600 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_292
timestamp 1607116009
transform 1 0 28244 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[113\]
timestamp 1607116009
transform 1 0 28612 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[260\]
timestamp 1607116009
transform 1 0 29348 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[27\]
timestamp 1607116009
transform 1 0 28888 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[374\]
timestamp 1607116009
transform 1 0 29624 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_302
timestamp 1607116009
transform 1 0 29164 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[167\]
timestamp 1607116009
transform 1 0 30176 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[385\]
timestamp 1607116009
transform 1 0 29900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[416\]
timestamp 1607116009
transform 1 0 30452 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[49\]
timestamp 1607116009
transform 1 0 30728 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[238\]
timestamp 1607116009
transform 1 0 31832 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_322
timestamp 1607116009
transform 1 0 31004 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_330
timestamp 1607116009
transform 1 0 31740 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[0\]
timestamp 1607116009
transform 1 0 32660 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[179\]
timestamp 1607116009
transform 1 0 33028 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[19\]
timestamp 1607116009
transform 1 0 32384 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_42
timestamp 1607116009
transform 1 0 32292 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_334
timestamp 1607116009
transform 1 0 32108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_343
timestamp 1607116009
transform 1 0 32936 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[332\]
timestamp 1607116009
transform 1 0 34316 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[389\]
timestamp 1607116009
transform 1 0 33304 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[77\]
timestamp 1607116009
transform 1 0 34040 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[80\]
timestamp 1607116009
transform 1 0 33580 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_353
timestamp 1607116009
transform 1 0 33856 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[206\]
timestamp 1607116009
transform 1 0 34684 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[41\]
timestamp 1607116009
transform 1 0 34960 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_361
timestamp 1607116009
transform 1 0 34592 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_368
timestamp 1607116009
transform 1 0 35236 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  insts\[8\]
timestamp 1607116009
transform 1 0 35880 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_374
timestamp 1607116009
transform 1 0 35788 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_378
timestamp 1607116009
transform 1 0 36156 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_43
timestamp 1607116009
transform 1 0 37904 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_390
timestamp 1607116009
transform 1 0 37260 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_396
timestamp 1607116009
transform 1 0 37812 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[45\]
timestamp 1607116009
transform 1 0 38456 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_398
timestamp 1607116009
transform 1 0 37996 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_402
timestamp 1607116009
transform 1 0 38364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_406
timestamp 1607116009
transform 1 0 38732 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_418
timestamp 1607116009
transform 1 0 39836 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[2\]
timestamp 1607116009
transform 1 0 40940 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_433
timestamp 1607116009
transform 1 0 41216 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[359\]
timestamp 1607116009
transform 1 0 41952 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_444
timestamp 1607116009
transform 1 0 42228 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_44
timestamp 1607116009
transform 1 0 43516 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_456
timestamp 1607116009
transform 1 0 43332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_459
timestamp 1607116009
transform 1 0 43608 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[94\]
timestamp 1607116009
transform 1 0 44528 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_467
timestamp 1607116009
transform 1 0 44344 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_472
timestamp 1607116009
transform 1 0 44804 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  insts\[79\]
timestamp 1607116009
transform 1 0 45172 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_479
timestamp 1607116009
transform 1 0 45448 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[434\]
timestamp 1607116009
transform 1 0 47104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_491
timestamp 1607116009
transform 1 0 46552 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_500
timestamp 1607116009
transform 1 0 47380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  insts\[78\]
timestamp 1607116009
transform 1 0 47840 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_504
timestamp 1607116009
transform 1 0 47748 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_508
timestamp 1607116009
transform 1 0 48116 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_45
timestamp 1607116009
transform 1 0 49128 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_516
timestamp 1607116009
transform 1 0 48852 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_520
timestamp 1607116009
transform 1 0 49220 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[81\]
timestamp 1607116009
transform 1 0 50324 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_535
timestamp 1607116009
transform 1 0 50600 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  insts\[443\]
timestamp 1607116009
transform 1 0 51152 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_544
timestamp 1607116009
transform 1 0 51428 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[376\]
timestamp 1607116009
transform 1 0 53268 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_556
timestamp 1607116009
transform 1 0 52532 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_567
timestamp 1607116009
transform 1 0 53544 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[418\]
timestamp 1607116009
transform 1 0 55384 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[427\]
timestamp 1607116009
transform 1 0 55660 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[54\]
timestamp 1607116009
transform 1 0 55108 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[57\]
timestamp 1607116009
transform 1 0 54832 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1607116009
transform 1 0 54740 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_579
timestamp 1607116009
transform 1 0 54648 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[226\]
timestamp 1607116009
transform 1 0 55936 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[250\]
timestamp 1607116009
transform 1 0 56212 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[322\]
timestamp 1607116009
transform 1 0 56488 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[396\]
timestamp 1607116009
transform 1 0 56764 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[99\]
timestamp 1607116009
transform 1 0 57040 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_608
timestamp 1607116009
transform 1 0 57316 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_616
timestamp 1607116009
transform 1 0 58052 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1607116009
transform -1 0 58604 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[70\]
timestamp 1607116009
transform 1 0 2484 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[90\]
timestamp 1607116009
transform 1 0 2208 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[95\]
timestamp 1607116009
transform 1 0 1932 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1607116009
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1607116009
transform 1 0 1656 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[16\]
timestamp 1607116009
transform 1 0 3588 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[193\]
timestamp 1607116009
transform 1 0 3312 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[292\]
timestamp 1607116009
transform 1 0 3036 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[312\]
timestamp 1607116009
transform 1 0 2760 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[133\]
timestamp 1607116009
transform 1 0 3864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[138\]
timestamp 1607116009
transform 1 0 4508 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[236\]
timestamp 1607116009
transform 1 0 4876 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1607116009
transform 1 0 4232 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_30
timestamp 1607116009
transform 1 0 4140 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_32
timestamp 1607116009
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_37
timestamp 1607116009
transform 1 0 4784 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[169\]
timestamp 1607116009
transform 1 0 5520 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[186\]
timestamp 1607116009
transform 1 0 5796 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[306\]
timestamp 1607116009
transform 1 0 5152 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[453\]
timestamp 1607116009
transform 1 0 6072 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_44
timestamp 1607116009
transform 1 0 5428 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[144\]
timestamp 1607116009
transform 1 0 6624 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[350\]
timestamp 1607116009
transform 1 0 6348 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[355\]
timestamp 1607116009
transform 1 0 7176 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1607116009
transform 1 0 7084 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_60
timestamp 1607116009
transform 1 0 6900 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[164\]
timestamp 1607116009
transform 1 0 8464 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[247\]
timestamp 1607116009
transform 1 0 7912 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[291\]
timestamp 1607116009
transform 1 0 8188 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[383\]
timestamp 1607116009
transform 1 0 7452 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_69
timestamp 1607116009
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[205\]
timestamp 1607116009
transform 1 0 8740 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[217\]
timestamp 1607116009
transform 1 0 9292 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[403\]
timestamp 1607116009
transform 1 0 9016 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_89
timestamp 1607116009
transform 1 0 9568 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[104\]
timestamp 1607116009
transform 1 0 10304 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[244\]
timestamp 1607116009
transform 1 0 10028 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[377\]
timestamp 1607116009
transform 1 0 10580 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[408\]
timestamp 1607116009
transform 1 0 9660 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1607116009
transform 1 0 9936 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[122\]
timestamp 1607116009
transform 1 0 11316 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[304\]
timestamp 1607116009
transform 1 0 11960 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[308\]
timestamp 1607116009
transform 1 0 11684 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[426\]
timestamp 1607116009
transform 1 0 10948 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_103
timestamp 1607116009
transform 1 0 10856 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_107
timestamp 1607116009
transform 1 0 11224 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1607116009
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[124\]
timestamp 1607116009
transform 1 0 12880 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[233\]
timestamp 1607116009
transform 1 0 12512 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[339\]
timestamp 1607116009
transform 1 0 12236 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1607116009
transform 1 0 12788 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_128
timestamp 1607116009
transform 1 0 13156 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[109\]
timestamp 1607116009
transform 1 0 14260 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[121\]
timestamp 1607116009
transform 1 0 13892 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[192\]
timestamp 1607116009
transform 1 0 13616 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[259\]
timestamp 1607116009
transform 1 0 13248 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_132
timestamp 1607116009
transform 1 0 13524 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_139
timestamp 1607116009
transform 1 0 14168 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[137\]
timestamp 1607116009
transform 1 0 14536 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[442\]
timestamp 1607116009
transform 1 0 15088 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[444\]
timestamp 1607116009
transform 1 0 15364 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[73\]
timestamp 1607116009
transform 1 0 14812 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[123\]
timestamp 1607116009
transform 1 0 16192 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[18\]
timestamp 1607116009
transform 1 0 15732 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[300\]
timestamp 1607116009
transform 1 0 16468 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1607116009
transform 1 0 15640 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_159
timestamp 1607116009
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[286\]
timestamp 1607116009
transform 1 0 17388 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[402\]
timestamp 1607116009
transform 1 0 17020 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[421\]
timestamp 1607116009
transform 1 0 16744 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[435\]
timestamp 1607116009
transform 1 0 17664 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_173
timestamp 1607116009
transform 1 0 17296 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[248\]
timestamp 1607116009
transform 1 0 18584 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[353\]
timestamp 1607116009
transform 1 0 18032 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[37\]
timestamp 1607116009
transform 1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1607116009
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_180
timestamp 1607116009
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_184
timestamp 1607116009
transform 1 0 18308 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[154\]
timestamp 1607116009
transform 1 0 20148 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[432\]
timestamp 1607116009
transform 1 0 19136 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[433\]
timestamp 1607116009
transform 1 0 19504 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[450\]
timestamp 1607116009
transform 1 0 19872 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_196
timestamp 1607116009
transform 1 0 19412 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_200
timestamp 1607116009
transform 1 0 19780 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[117\]
timestamp 1607116009
transform 1 0 20516 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[131\]
timestamp 1607116009
transform 1 0 21436 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[148\]
timestamp 1607116009
transform 1 0 20792 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[53\]
timestamp 1607116009
transform 1 0 21068 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1607116009
transform 1 0 21344 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_207
timestamp 1607116009
transform 1 0 20424 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[107\]
timestamp 1607116009
transform 1 0 21804 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[347\]
timestamp 1607116009
transform 1 0 22080 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[395\]
timestamp 1607116009
transform 1 0 22356 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[58\]
timestamp 1607116009
transform 1 0 22632 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_221
timestamp 1607116009
transform 1 0 21712 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[74\]
timestamp 1607116009
transform 1 0 22908 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[84\]
timestamp 1607116009
transform 1 0 23184 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[87\]
timestamp 1607116009
transform 1 0 23552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_240
timestamp 1607116009
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[454\]
timestamp 1607116009
transform 1 0 24288 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[98\]
timestamp 1607116009
transform 1 0 23828 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1607116009
transform 1 0 24196 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_247
timestamp 1607116009
transform 1 0 24104 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_252
timestamp 1607116009
transform 1 0 24564 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[445\]
timestamp 1607116009
transform 1 0 25576 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_260
timestamp 1607116009
transform 1 0 25300 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_266
timestamp 1607116009
transform 1 0 25852 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1607116009
transform 1 0 27048 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_278
timestamp 1607116009
transform 1 0 26956 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_280
timestamp 1607116009
transform 1 0 27140 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[366\]
timestamp 1607116009
transform 1 0 28152 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[398\]
timestamp 1607116009
transform 1 0 28428 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_288
timestamp 1607116009
transform 1 0 27876 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[364\]
timestamp 1607116009
transform 1 0 28704 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_300
timestamp 1607116009
transform 1 0 28980 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_308
timestamp 1607116009
transform 1 0 29716 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[340\]
timestamp 1607116009
transform 1 0 30636 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1607116009
transform 1 0 29900 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_311
timestamp 1607116009
transform 1 0 29992 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_317
timestamp 1607116009
transform 1 0 30544 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[431\]
timestamp 1607116009
transform 1 0 31832 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[5\]
timestamp 1607116009
transform 1 0 31556 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_321
timestamp 1607116009
transform 1 0 30912 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_327
timestamp 1607116009
transform 1 0 31464 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[152\]
timestamp 1607116009
transform 1 0 32108 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[188\]
timestamp 1607116009
transform 1 0 32844 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[309\]
timestamp 1607116009
transform 1 0 32384 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[328\]
timestamp 1607116009
transform 1 0 33120 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1607116009
transform 1 0 32752 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_340
timestamp 1607116009
transform 1 0 32660 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[338\]
timestamp 1607116009
transform 1 0 34224 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[358\]
timestamp 1607116009
transform 1 0 33396 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[430\]
timestamp 1607116009
transform 1 0 33672 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_354
timestamp 1607116009
transform 1 0 33948 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[163\]
timestamp 1607116009
transform 1 0 34960 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[210\]
timestamp 1607116009
transform 1 0 34500 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[273\]
timestamp 1607116009
transform 1 0 35236 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1607116009
transform 1 0 35604 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_363
timestamp 1607116009
transform 1 0 34776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_371
timestamp 1607116009
transform 1 0 35512 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[11\]
timestamp 1607116009
transform 1 0 36248 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[127\]
timestamp 1607116009
transform 1 0 35696 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[380\]
timestamp 1607116009
transform 1 0 36524 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[409\]
timestamp 1607116009
transform 1 0 35972 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_385
timestamp 1607116009
transform 1 0 36800 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[140\]
timestamp 1607116009
transform 1 0 36892 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[151\]
timestamp 1607116009
transform 1 0 37628 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[165\]
timestamp 1607116009
transform 1 0 37168 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[230\]
timestamp 1607116009
transform 1 0 37904 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_392
timestamp 1607116009
transform 1 0 37444 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[130\]
timestamp 1607116009
transform 1 0 38548 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[288\]
timestamp 1607116009
transform 1 0 38824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[290\]
timestamp 1607116009
transform 1 0 38180 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[333\]
timestamp 1607116009
transform 1 0 39100 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1607116009
transform 1 0 38456 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[189\]
timestamp 1607116009
transform 1 0 39376 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[196\]
timestamp 1607116009
transform 1 0 40020 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[24\]
timestamp 1607116009
transform 1 0 39652 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_419
timestamp 1607116009
transform 1 0 39928 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_423
timestamp 1607116009
transform 1 0 40296 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[174\]
timestamp 1607116009
transform 1 0 40756 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[241\]
timestamp 1607116009
transform 1 0 40388 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[275\]
timestamp 1607116009
transform 1 0 41032 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1607116009
transform 1 0 41308 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_427
timestamp 1607116009
transform 1 0 40664 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_435
timestamp 1607116009
transform 1 0 41400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[135\]
timestamp 1607116009
transform 1 0 41584 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[145\]
timestamp 1607116009
transform 1 0 42228 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[162\]
timestamp 1607116009
transform 1 0 42596 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[274\]
timestamp 1607116009
transform 1 0 41860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_443
timestamp 1607116009
transform 1 0 42136 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1607116009
transform 1 0 42504 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[224\]
timestamp 1607116009
transform 1 0 42872 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[337\]
timestamp 1607116009
transform 1 0 43608 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[354\]
timestamp 1607116009
transform 1 0 43884 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[76\]
timestamp 1607116009
transform 1 0 43148 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_457
timestamp 1607116009
transform 1 0 43424 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[126\]
timestamp 1607116009
transform 1 0 44804 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[256\]
timestamp 1607116009
transform 1 0 44252 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[387\]
timestamp 1607116009
transform 1 0 44528 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1607116009
transform 1 0 44160 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[118\]
timestamp 1607116009
transform 1 0 45540 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[229\]
timestamp 1607116009
transform 1 0 46000 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[441\]
timestamp 1607116009
transform 1 0 45264 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_475
timestamp 1607116009
transform 1 0 45080 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_483
timestamp 1607116009
transform 1 0 45816 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[252\]
timestamp 1607116009
transform 1 0 46552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[269\]
timestamp 1607116009
transform 1 0 47288 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[393\]
timestamp 1607116009
transform 1 0 46276 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1607116009
transform 1 0 47012 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_494
timestamp 1607116009
transform 1 0 46828 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_497
timestamp 1607116009
transform 1 0 47104 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[257\]
timestamp 1607116009
transform 1 0 48024 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[352\]
timestamp 1607116009
transform 1 0 47564 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[52\]
timestamp 1607116009
transform 1 0 48300 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_505
timestamp 1607116009
transform 1 0 47840 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_513
timestamp 1607116009
transform 1 0 48576 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[356\]
timestamp 1607116009
transform 1 0 49312 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[370\]
timestamp 1607116009
transform 1 0 48668 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[60\]
timestamp 1607116009
transform 1 0 49588 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[75\]
timestamp 1607116009
transform 1 0 48944 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_520
timestamp 1607116009
transform 1 0 49220 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[111\]
timestamp 1607116009
transform 1 0 50692 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[227\]
timestamp 1607116009
transform 1 0 49956 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[243\]
timestamp 1607116009
transform 1 0 50232 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[32\]
timestamp 1607116009
transform 1 0 50968 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1607116009
transform 1 0 49864 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_534
timestamp 1607116009
transform 1 0 50508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[155\]
timestamp 1607116009
transform 1 0 51336 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[183\]
timestamp 1607116009
transform 1 0 51704 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[316\]
timestamp 1607116009
transform 1 0 51980 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_542
timestamp 1607116009
transform 1 0 51244 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_546
timestamp 1607116009
transform 1 0 51612 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[161\]
timestamp 1607116009
transform 1 0 52808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[298\]
timestamp 1607116009
transform 1 0 53084 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[88\]
timestamp 1607116009
transform 1 0 52348 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1607116009
transform 1 0 52716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_553
timestamp 1607116009
transform 1 0 52256 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_557
timestamp 1607116009
transform 1 0 52624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[128\]
timestamp 1607116009
transform 1 0 53912 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[134\]
timestamp 1607116009
transform 1 0 54188 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[35\]
timestamp 1607116009
transform 1 0 53544 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[438\]
timestamp 1607116009
transform 1 0 54464 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_565
timestamp 1607116009
transform 1 0 53360 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_570
timestamp 1607116009
transform 1 0 53820 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[173\]
timestamp 1607116009
transform 1 0 55108 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[218\]
timestamp 1607116009
transform 1 0 54740 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[271\]
timestamp 1607116009
transform 1 0 55660 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1607116009
transform 1 0 55568 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_583
timestamp 1607116009
transform 1 0 55016 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_587
timestamp 1607116009
transform 1 0 55384 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[136\]
timestamp 1607116009
transform 1 0 55936 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[141\]
timestamp 1607116009
transform 1 0 56212 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[147\]
timestamp 1607116009
transform 1 0 56488 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[242\]
timestamp 1607116009
transform 1 0 56764 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[336\]
timestamp 1607116009
transform 1 0 57040 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[404\]
timestamp 1607116009
transform 1 0 57316 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[425\]
timestamp 1607116009
transform 1 0 57592 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_614
timestamp 1607116009
transform 1 0 57868 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1607116009
transform -1 0 58604 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_618
timestamp 1607116009
transform 1 0 58236 0 1 2720
box -38 -48 130 592
<< labels >>
rlabel metal2 s 32954 3800 33010 4600 6 HI[0]
port 0 nsew signal tristate
rlabel metal3 s 59200 1912 60000 2032 6 HI[100]
port 1 nsew signal tristate
rlabel metal2 s 28906 3800 28962 4600 6 HI[101]
port 2 nsew signal tristate
rlabel metal2 s 35714 0 35770 800 6 HI[102]
port 3 nsew signal tristate
rlabel metal2 s 25410 0 25466 800 6 HI[103]
port 4 nsew signal tristate
rlabel metal2 s 9402 3800 9458 4600 6 HI[104]
port 5 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 HI[105]
port 6 nsew signal tristate
rlabel metal2 s 9954 0 10010 800 6 HI[106]
port 7 nsew signal tristate
rlabel metal2 s 20442 3800 20498 4600 6 HI[107]
port 8 nsew signal tristate
rlabel metal2 s 42706 0 42762 800 6 HI[108]
port 9 nsew signal tristate
rlabel metal2 s 13082 3800 13138 4600 6 HI[109]
port 10 nsew signal tristate
rlabel metal2 s 54850 0 54906 800 6 HI[10]
port 11 nsew signal tristate
rlabel metal2 s 3698 0 3754 800 6 HI[110]
port 12 nsew signal tristate
rlabel metal2 s 51722 3800 51778 4600 6 HI[111]
port 13 nsew signal tristate
rlabel metal2 s 9218 0 9274 800 6 HI[112]
port 14 nsew signal tristate
rlabel metal2 s 28170 3800 28226 4600 6 HI[113]
port 15 nsew signal tristate
rlabel metal2 s 46386 0 46442 800 6 HI[114]
port 16 nsew signal tristate
rlabel metal2 s 12898 0 12954 800 6 HI[115]
port 17 nsew signal tristate
rlabel metal2 s 5538 0 5594 800 6 HI[116]
port 18 nsew signal tristate
rlabel metal2 s 18970 3800 19026 4600 6 HI[117]
port 19 nsew signal tristate
rlabel metal2 s 46938 3800 46994 4600 6 HI[118]
port 20 nsew signal tristate
rlabel metal2 s 10874 0 10930 800 6 HI[119]
port 21 nsew signal tristate
rlabel metal2 s 38290 3800 38346 4600 6 HI[11]
port 22 nsew signal tristate
rlabel metal2 s 41786 0 41842 800 6 HI[120]
port 23 nsew signal tristate
rlabel metal2 s 12714 3800 12770 4600 6 HI[121]
port 24 nsew signal tristate
rlabel metal2 s 10322 3800 10378 4600 6 HI[122]
port 25 nsew signal tristate
rlabel metal2 s 14922 3800 14978 4600 6 HI[123]
port 26 nsew signal tristate
rlabel metal2 s 11794 3800 11850 4600 6 HI[124]
port 27 nsew signal tristate
rlabel metal2 s 22282 0 22338 800 6 HI[125]
port 28 nsew signal tristate
rlabel metal2 s 46202 3800 46258 4600 6 HI[126]
port 29 nsew signal tristate
rlabel metal2 s 37738 3800 37794 4600 6 HI[127]
port 30 nsew signal tristate
rlabel metal2 s 54482 3800 54538 4600 6 HI[128]
port 31 nsew signal tristate
rlabel metal2 s 18050 0 18106 800 6 HI[129]
port 32 nsew signal tristate
rlabel metal2 s 7378 0 7434 800 6 HI[12]
port 33 nsew signal tristate
rlabel metal2 s 40130 3800 40186 4600 6 HI[130]
port 34 nsew signal tristate
rlabel metal2 s 19706 3800 19762 4600 6 HI[131]
port 35 nsew signal tristate
rlabel metal2 s 33874 0 33930 800 6 HI[132]
port 36 nsew signal tristate
rlabel metal2 s 3698 3800 3754 4600 6 HI[133]
port 37 nsew signal tristate
rlabel metal2 s 54666 3800 54722 4600 6 HI[134]
port 38 nsew signal tristate
rlabel metal2 s 43258 3800 43314 4600 6 HI[135]
port 39 nsew signal tristate
rlabel metal2 s 58346 3800 58402 4600 6 HI[136]
port 40 nsew signal tristate
rlabel metal2 s 13266 3800 13322 4600 6 HI[137]
port 41 nsew signal tristate
rlabel metal2 s 4250 3800 4306 4600 6 HI[138]
port 42 nsew signal tristate
rlabel metal2 s 9034 0 9090 800 6 HI[139]
port 43 nsew signal tristate
rlabel metal2 s 50434 0 50490 800 6 HI[13]
port 44 nsew signal tristate
rlabel metal2 s 38842 3800 38898 4600 6 HI[140]
port 45 nsew signal tristate
rlabel metal2 s 58898 3800 58954 4600 6 HI[141]
port 46 nsew signal tristate
rlabel metal2 s 34794 0 34850 800 6 HI[142]
port 47 nsew signal tristate
rlabel metal2 s 6826 0 6882 800 6 HI[143]
port 48 nsew signal tristate
rlabel metal2 s 6090 3800 6146 4600 6 HI[144]
port 49 nsew signal tristate
rlabel metal2 s 43810 3800 43866 4600 6 HI[145]
port 50 nsew signal tristate
rlabel metal2 s 26330 3800 26386 4600 6 HI[146]
port 51 nsew signal tristate
rlabel metal2 s 59266 3800 59322 4600 6 HI[147]
port 52 nsew signal tristate
rlabel metal2 s 19154 3800 19210 4600 6 HI[148]
port 53 nsew signal tristate
rlabel metal2 s 11426 0 11482 800 6 HI[149]
port 54 nsew signal tristate
rlabel metal2 s 36082 0 36138 800 6 HI[14]
port 55 nsew signal tristate
rlabel metal2 s 28906 0 28962 800 6 HI[150]
port 56 nsew signal tristate
rlabel metal2 s 39578 3800 39634 4600 6 HI[151]
port 57 nsew signal tristate
rlabel metal2 s 34794 3800 34850 4600 6 HI[152]
port 58 nsew signal tristate
rlabel metal2 s 43258 0 43314 800 6 HI[153]
port 59 nsew signal tristate
rlabel metal2 s 18602 3800 18658 4600 6 HI[154]
port 60 nsew signal tristate
rlabel metal2 s 52274 3800 52330 4600 6 HI[155]
port 61 nsew signal tristate
rlabel metal2 s 26146 0 26202 800 6 HI[156]
port 62 nsew signal tristate
rlabel metal2 s 30010 0 30066 800 6 HI[157]
port 63 nsew signal tristate
rlabel metal2 s 56506 0 56562 800 6 HI[158]
port 64 nsew signal tristate
rlabel metal2 s 7562 0 7618 800 6 HI[159]
port 65 nsew signal tristate
rlabel metal2 s 25778 0 25834 800 6 HI[15]
port 66 nsew signal tristate
rlabel metal2 s 14186 0 14242 800 6 HI[160]
port 67 nsew signal tristate
rlabel metal2 s 53378 3800 53434 4600 6 HI[161]
port 68 nsew signal tristate
rlabel metal2 s 44178 3800 44234 4600 6 HI[162]
port 69 nsew signal tristate
rlabel metal2 s 37002 3800 37058 4600 6 HI[163]
port 70 nsew signal tristate
rlabel metal2 s 7746 3800 7802 4600 6 HI[164]
port 71 nsew signal tristate
rlabel metal2 s 39026 3800 39082 4600 6 HI[165]
port 72 nsew signal tristate
rlabel metal2 s 23018 0 23074 800 6 HI[166]
port 73 nsew signal tristate
rlabel metal2 s 30562 3800 30618 4600 6 HI[167]
port 74 nsew signal tristate
rlabel metal2 s 9770 0 9826 800 6 HI[168]
port 75 nsew signal tristate
rlabel metal2 s 5170 3800 5226 4600 6 HI[169]
port 76 nsew signal tristate
rlabel metal2 s 2962 3800 3018 4600 6 HI[16]
port 77 nsew signal tristate
rlabel metal2 s 12162 0 12218 800 6 HI[170]
port 78 nsew signal tristate
rlabel metal2 s 33322 0 33378 800 6 HI[171]
port 79 nsew signal tristate
rlabel metal2 s 34978 0 35034 800 6 HI[172]
port 80 nsew signal tristate
rlabel metal2 s 55586 3800 55642 4600 6 HI[173]
port 81 nsew signal tristate
rlabel metal2 s 42522 3800 42578 4600 6 HI[174]
port 82 nsew signal tristate
rlabel metal2 s 47490 0 47546 800 6 HI[175]
port 83 nsew signal tristate
rlabel metal2 s 938 0 994 800 6 HI[176]
port 84 nsew signal tristate
rlabel metal2 s 4986 0 5042 800 6 HI[177]
port 85 nsew signal tristate
rlabel metal2 s 21546 3800 21602 4600 6 HI[178]
port 86 nsew signal tristate
rlabel metal2 s 33138 3800 33194 4600 6 HI[179]
port 87 nsew signal tristate
rlabel metal2 s 27066 0 27122 800 6 HI[17]
port 88 nsew signal tristate
rlabel metal2 s 5722 0 5778 800 6 HI[180]
port 89 nsew signal tristate
rlabel metal2 s 11610 0 11666 800 6 HI[181]
port 90 nsew signal tristate
rlabel metal2 s 39026 0 39082 800 6 HI[182]
port 91 nsew signal tristate
rlabel metal2 s 52642 3800 52698 4600 6 HI[183]
port 92 nsew signal tristate
rlabel metal2 s 24674 3800 24730 4600 6 HI[184]
port 93 nsew signal tristate
rlabel metal2 s 9586 0 9642 800 6 HI[185]
port 94 nsew signal tristate
rlabel metal2 s 5354 3800 5410 4600 6 HI[186]
port 95 nsew signal tristate
rlabel metal2 s 10506 0 10562 800 6 HI[187]
port 96 nsew signal tristate
rlabel metal2 s 35530 3800 35586 4600 6 HI[188]
port 97 nsew signal tristate
rlabel metal2 s 41234 3800 41290 4600 6 HI[189]
port 98 nsew signal tristate
rlabel metal2 s 14370 3800 14426 4600 6 HI[18]
port 99 nsew signal tristate
rlabel metal2 s 53010 0 53066 800 6 HI[190]
port 100 nsew signal tristate
rlabel metal2 s 22650 3800 22706 4600 6 HI[191]
port 101 nsew signal tristate
rlabel metal2 s 12530 3800 12586 4600 6 HI[192]
port 102 nsew signal tristate
rlabel metal2 s 1674 3800 1730 4600 6 HI[193]
port 103 nsew signal tristate
rlabel metal2 s 54666 0 54722 800 6 HI[194]
port 104 nsew signal tristate
rlabel metal2 s 38658 0 38714 800 6 HI[195]
port 105 nsew signal tristate
rlabel metal2 s 41786 3800 41842 4600 6 HI[196]
port 106 nsew signal tristate
rlabel metal2 s 23386 3800 23442 4600 6 HI[197]
port 107 nsew signal tristate
rlabel metal2 s 58898 0 58954 800 6 HI[198]
port 108 nsew signal tristate
rlabel metal2 s 29458 0 29514 800 6 HI[199]
port 109 nsew signal tristate
rlabel metal2 s 31666 3800 31722 4600 6 HI[19]
port 110 nsew signal tristate
rlabel metal2 s 12346 0 12402 800 6 HI[1]
port 111 nsew signal tristate
rlabel metal2 s 26698 0 26754 800 6 HI[200]
port 112 nsew signal tristate
rlabel metal3 s 0 1912 800 2032 6 HI[201]
port 113 nsew signal tristate
rlabel metal2 s 23386 0 23442 800 6 HI[202]
port 114 nsew signal tristate
rlabel metal2 s 52274 0 52330 800 6 HI[203]
port 115 nsew signal tristate
rlabel metal2 s 47122 0 47178 800 6 HI[204]
port 116 nsew signal tristate
rlabel metal2 s 7930 3800 7986 4600 6 HI[205]
port 117 nsew signal tristate
rlabel metal2 s 34058 3800 34114 4600 6 HI[206]
port 118 nsew signal tristate
rlabel metal2 s 24122 3800 24178 4600 6 HI[207]
port 119 nsew signal tristate
rlabel metal2 s 37370 0 37426 800 6 HI[208]
port 120 nsew signal tristate
rlabel metal2 s 45282 0 45338 800 6 HI[209]
port 121 nsew signal tristate
rlabel metal2 s 56690 0 56746 800 6 HI[20]
port 122 nsew signal tristate
rlabel metal2 s 36634 3800 36690 4600 6 HI[210]
port 123 nsew signal tristate
rlabel metal2 s 19522 0 19578 800 6 HI[211]
port 124 nsew signal tristate
rlabel metal2 s 17498 0 17554 800 6 HI[212]
port 125 nsew signal tristate
rlabel metal2 s 1306 0 1362 800 6 HI[213]
port 126 nsew signal tristate
rlabel metal2 s 27986 0 28042 800 6 HI[214]
port 127 nsew signal tristate
rlabel metal2 s 39762 0 39818 800 6 HI[215]
port 128 nsew signal tristate
rlabel metal2 s 42338 0 42394 800 6 HI[216]
port 129 nsew signal tristate
rlabel metal2 s 8482 3800 8538 4600 6 HI[217]
port 130 nsew signal tristate
rlabel metal2 s 55218 3800 55274 4600 6 HI[218]
port 131 nsew signal tristate
rlabel metal2 s 7930 0 7986 800 6 HI[219]
port 132 nsew signal tristate
rlabel metal2 s 27618 3800 27674 4600 6 HI[21]
port 133 nsew signal tristate
rlabel metal2 s 30746 0 30802 800 6 HI[220]
port 134 nsew signal tristate
rlabel metal2 s 3330 0 3386 800 6 HI[221]
port 135 nsew signal tristate
rlabel metal2 s 40498 0 40554 800 6 HI[222]
port 136 nsew signal tristate
rlabel metal3 s 0 2184 800 2304 6 HI[223]
port 137 nsew signal tristate
rlabel metal2 s 44362 3800 44418 4600 6 HI[224]
port 138 nsew signal tristate
rlabel metal2 s 754 3800 810 4600 6 HI[225]
port 139 nsew signal tristate
rlabel metal3 s 59200 3000 60000 3120 6 HI[226]
port 140 nsew signal tristate
rlabel metal2 s 50802 3800 50858 4600 6 HI[227]
port 141 nsew signal tristate
rlabel metal2 s 45834 0 45890 800 6 HI[228]
port 142 nsew signal tristate
rlabel metal2 s 47306 3800 47362 4600 6 HI[229]
port 143 nsew signal tristate
rlabel metal2 s 20442 0 20498 800 6 HI[22]
port 144 nsew signal tristate
rlabel metal2 s 39394 3800 39450 4600 6 HI[230]
port 145 nsew signal tristate
rlabel metal2 s 12714 0 12770 800 6 HI[231]
port 146 nsew signal tristate
rlabel metal2 s 11978 0 12034 800 6 HI[232]
port 147 nsew signal tristate
rlabel metal2 s 11426 3800 11482 4600 6 HI[233]
port 148 nsew signal tristate
rlabel metal2 s 49882 0 49938 800 6 HI[234]
port 149 nsew signal tristate
rlabel metal2 s 3882 0 3938 800 6 HI[235]
port 150 nsew signal tristate
rlabel metal2 s 4618 3800 4674 4600 6 HI[236]
port 151 nsew signal tristate
rlabel metal2 s 43442 0 43498 800 6 HI[237]
port 152 nsew signal tristate
rlabel metal2 s 31298 3800 31354 4600 6 HI[238]
port 153 nsew signal tristate
rlabel metal2 s 54298 0 54354 800 6 HI[239]
port 154 nsew signal tristate
rlabel metal2 s 31298 0 31354 800 6 HI[23]
port 155 nsew signal tristate
rlabel metal2 s 4434 0 4490 800 6 HI[240]
port 156 nsew signal tristate
rlabel metal2 s 42154 3800 42210 4600 6 HI[241]
port 157 nsew signal tristate
rlabel metal2 s 56322 3800 56378 4600 6 HI[242]
port 158 nsew signal tristate
rlabel metal2 s 50986 3800 51042 4600 6 HI[243]
port 159 nsew signal tristate
rlabel metal2 s 9034 3800 9090 4600 6 HI[244]
port 160 nsew signal tristate
rlabel metal2 s 17130 0 17186 800 6 HI[245]
port 161 nsew signal tristate
rlabel metal2 s 54114 0 54170 800 6 HI[246]
port 162 nsew signal tristate
rlabel metal2 s 7194 3800 7250 4600 6 HI[247]
port 163 nsew signal tristate
rlabel metal2 s 16946 3800 17002 4600 6 HI[248]
port 164 nsew signal tristate
rlabel metal2 s 14738 0 14794 800 6 HI[249]
port 165 nsew signal tristate
rlabel metal2 s 41418 3800 41474 4600 6 HI[24]
port 166 nsew signal tristate
rlabel metal3 s 59200 3544 60000 3664 6 HI[250]
port 167 nsew signal tristate
rlabel metal2 s 16578 0 16634 800 6 HI[251]
port 168 nsew signal tristate
rlabel metal2 s 47858 3800 47914 4600 6 HI[252]
port 169 nsew signal tristate
rlabel metal2 s 25594 3800 25650 4600 6 HI[253]
port 170 nsew signal tristate
rlabel metal2 s 27250 0 27306 800 6 HI[254]
port 171 nsew signal tristate
rlabel metal2 s 48778 0 48834 800 6 HI[255]
port 172 nsew signal tristate
rlabel metal2 s 45466 3800 45522 4600 6 HI[256]
port 173 nsew signal tristate
rlabel metal2 s 49330 3800 49386 4600 6 HI[257]
port 174 nsew signal tristate
rlabel metal2 s 4250 0 4306 800 6 HI[258]
port 175 nsew signal tristate
rlabel metal2 s 12162 3800 12218 4600 6 HI[259]
port 176 nsew signal tristate
rlabel metal2 s 21730 3800 21786 4600 6 HI[25]
port 177 nsew signal tristate
rlabel metal2 s 29826 3800 29882 4600 6 HI[260]
port 178 nsew signal tristate
rlabel metal2 s 51170 0 51226 800 6 HI[261]
port 179 nsew signal tristate
rlabel metal2 s 53378 0 53434 800 6 HI[262]
port 180 nsew signal tristate
rlabel metal2 s 22282 3800 22338 4600 6 HI[263]
port 181 nsew signal tristate
rlabel metal2 s 52458 0 52514 800 6 HI[264]
port 182 nsew signal tristate
rlabel metal2 s 15106 0 15162 800 6 HI[265]
port 183 nsew signal tristate
rlabel metal2 s 37922 0 37978 800 6 HI[266]
port 184 nsew signal tristate
rlabel metal2 s 25962 3800 26018 4600 6 HI[267]
port 185 nsew signal tristate
rlabel metal2 s 570 0 626 800 6 HI[268]
port 186 nsew signal tristate
rlabel metal2 s 48594 3800 48650 4600 6 HI[269]
port 187 nsew signal tristate
rlabel metal2 s 6090 0 6146 800 6 HI[26]
port 188 nsew signal tristate
rlabel metal2 s 3146 0 3202 800 6 HI[270]
port 189 nsew signal tristate
rlabel metal2 s 56874 3800 56930 4600 6 HI[271]
port 190 nsew signal tristate
rlabel metal2 s 27434 3800 27490 4600 6 HI[272]
port 191 nsew signal tristate
rlabel metal2 s 37186 3800 37242 4600 6 HI[273]
port 192 nsew signal tristate
rlabel metal2 s 43074 3800 43130 4600 6 HI[274]
port 193 nsew signal tristate
rlabel metal2 s 41970 3800 42026 4600 6 HI[275]
port 194 nsew signal tristate
rlabel metal2 s 40866 0 40922 800 6 HI[276]
port 195 nsew signal tristate
rlabel metal2 s 45098 0 45154 800 6 HI[277]
port 196 nsew signal tristate
rlabel metal2 s 34242 0 34298 800 6 HI[278]
port 197 nsew signal tristate
rlabel metal2 s 55402 0 55458 800 6 HI[279]
port 198 nsew signal tristate
rlabel metal2 s 28354 3800 28410 4600 6 HI[27]
port 199 nsew signal tristate
rlabel metal2 s 48226 0 48282 800 6 HI[280]
port 200 nsew signal tristate
rlabel metal2 s 1306 3800 1362 4600 6 HI[281]
port 201 nsew signal tristate
rlabel metal2 s 27066 3800 27122 4600 6 HI[282]
port 202 nsew signal tristate
rlabel metal2 s 36818 0 36874 800 6 HI[283]
port 203 nsew signal tristate
rlabel metal2 s 30378 0 30434 800 6 HI[284]
port 204 nsew signal tristate
rlabel metal3 s 59200 2184 60000 2304 6 HI[285]
port 205 nsew signal tristate
rlabel metal2 s 16026 3800 16082 4600 6 HI[286]
port 206 nsew signal tristate
rlabel metal2 s 25226 3800 25282 4600 6 HI[287]
port 207 nsew signal tristate
rlabel metal2 s 40682 3800 40738 4600 6 HI[288]
port 208 nsew signal tristate
rlabel metal2 s 22098 3800 22154 4600 6 HI[289]
port 209 nsew signal tristate
rlabel metal2 s 38106 0 38162 800 6 HI[28]
port 210 nsew signal tristate
rlabel metal2 s 39762 3800 39818 4600 6 HI[290]
port 211 nsew signal tristate
rlabel metal2 s 7010 3800 7066 4600 6 HI[291]
port 212 nsew signal tristate
rlabel metal2 s 2410 3800 2466 4600 6 HI[292]
port 213 nsew signal tristate
rlabel metal2 s 18602 0 18658 800 6 HI[293]
port 214 nsew signal tristate
rlabel metal2 s 58346 0 58402 800 6 HI[294]
port 215 nsew signal tristate
rlabel metal2 s 50066 0 50122 800 6 HI[295]
port 216 nsew signal tristate
rlabel metal2 s 40314 0 40370 800 6 HI[296]
port 217 nsew signal tristate
rlabel metal2 s 42154 0 42210 800 6 HI[297]
port 218 nsew signal tristate
rlabel metal2 s 53562 3800 53618 4600 6 HI[298]
port 219 nsew signal tristate
rlabel metal2 s 37554 0 37610 800 6 HI[299]
port 220 nsew signal tristate
rlabel metal2 s 46202 0 46258 800 6 HI[29]
port 221 nsew signal tristate
rlabel metal2 s 42706 3800 42762 4600 6 HI[2]
port 222 nsew signal tristate
rlabel metal2 s 14554 3800 14610 4600 6 HI[300]
port 223 nsew signal tristate
rlabel metal2 s 2594 0 2650 800 6 HI[301]
port 224 nsew signal tristate
rlabel metal2 s 27618 0 27674 800 6 HI[302]
port 225 nsew signal tristate
rlabel metal2 s 39578 0 39634 800 6 HI[303]
port 226 nsew signal tristate
rlabel metal2 s 10874 3800 10930 4600 6 HI[304]
port 227 nsew signal tristate
rlabel metal2 s 37186 0 37242 800 6 HI[305]
port 228 nsew signal tristate
rlabel metal2 s 4802 3800 4858 4600 6 HI[306]
port 229 nsew signal tristate
rlabel metal2 s 44546 0 44602 800 6 HI[307]
port 230 nsew signal tristate
rlabel metal2 s 10690 3800 10746 4600 6 HI[308]
port 231 nsew signal tristate
rlabel metal2 s 32770 3800 32826 4600 6 HI[309]
port 232 nsew signal tristate
rlabel metal2 s 41602 0 41658 800 6 HI[30]
port 233 nsew signal tristate
rlabel metal2 s 8114 0 8170 800 6 HI[310]
port 234 nsew signal tristate
rlabel metal2 s 18970 0 19026 800 6 HI[311]
port 235 nsew signal tristate
rlabel metal2 s 2226 3800 2282 4600 6 HI[312]
port 236 nsew signal tristate
rlabel metal2 s 53746 0 53802 800 6 HI[313]
port 237 nsew signal tristate
rlabel metal2 s 11058 0 11114 800 6 HI[314]
port 238 nsew signal tristate
rlabel metal2 s 32770 0 32826 800 6 HI[315]
port 239 nsew signal tristate
rlabel metal2 s 52826 3800 52882 4600 6 HI[316]
port 240 nsew signal tristate
rlabel metal2 s 8666 0 8722 800 6 HI[317]
port 241 nsew signal tristate
rlabel metal2 s 22834 0 22890 800 6 HI[318]
port 242 nsew signal tristate
rlabel metal2 s 42890 0 42946 800 6 HI[319]
port 243 nsew signal tristate
rlabel metal2 s 47674 0 47730 800 6 HI[31]
port 244 nsew signal tristate
rlabel metal2 s 6274 0 6330 800 6 HI[320]
port 245 nsew signal tristate
rlabel metal2 s 2778 0 2834 800 6 HI[321]
port 246 nsew signal tristate
rlabel metal2 s 57610 3800 57666 4600 6 HI[322]
port 247 nsew signal tristate
rlabel metal2 s 6642 0 6698 800 6 HI[323]
port 248 nsew signal tristate
rlabel metal2 s 15290 0 15346 800 6 HI[324]
port 249 nsew signal tristate
rlabel metal2 s 23754 3800 23810 4600 6 HI[325]
port 250 nsew signal tristate
rlabel metal2 s 32034 0 32090 800 6 HI[326]
port 251 nsew signal tristate
rlabel metal2 s 23754 0 23810 800 6 HI[327]
port 252 nsew signal tristate
rlabel metal2 s 35898 3800 35954 4600 6 HI[328]
port 253 nsew signal tristate
rlabel metal2 s 24674 0 24730 800 6 HI[329]
port 254 nsew signal tristate
rlabel metal2 s 51538 3800 51594 4600 6 HI[32]
port 255 nsew signal tristate
rlabel metal2 s 28538 0 28594 800 6 HI[330]
port 256 nsew signal tristate
rlabel metal2 s 14002 0 14058 800 6 HI[331]
port 257 nsew signal tristate
rlabel metal2 s 33690 3800 33746 4600 6 HI[332]
port 258 nsew signal tristate
rlabel metal2 s 40866 3800 40922 4600 6 HI[333]
port 259 nsew signal tristate
rlabel metal2 s 32586 0 32642 800 6 HI[334]
port 260 nsew signal tristate
rlabel metal2 s 58530 0 58586 800 6 HI[335]
port 261 nsew signal tristate
rlabel metal2 s 57978 3800 58034 4600 6 HI[336]
port 262 nsew signal tristate
rlabel metal2 s 45098 3800 45154 4600 6 HI[337]
port 263 nsew signal tristate
rlabel metal2 s 36450 3800 36506 4600 6 HI[338]
port 264 nsew signal tristate
rlabel metal2 s 11242 3800 11298 4600 6 HI[339]
port 265 nsew signal tristate
rlabel metal3 s 0 3000 800 3120 6 HI[33]
port 266 nsew signal tristate
rlabel metal2 s 32402 3800 32458 4600 6 HI[340]
port 267 nsew signal tristate
rlabel metal2 s 15658 0 15714 800 6 HI[341]
port 268 nsew signal tristate
rlabel metal2 s 25042 3800 25098 4600 6 HI[342]
port 269 nsew signal tristate
rlabel metal2 s 53562 0 53618 800 6 HI[343]
port 270 nsew signal tristate
rlabel metal2 s 23570 0 23626 800 6 HI[344]
port 271 nsew signal tristate
rlabel metal2 s 39946 0 40002 800 6 HI[345]
port 272 nsew signal tristate
rlabel metal2 s 4802 0 4858 800 6 HI[346]
port 273 nsew signal tristate
rlabel metal2 s 19890 3800 19946 4600 6 HI[347]
port 274 nsew signal tristate
rlabel metal2 s 23938 3800 23994 4600 6 HI[348]
port 275 nsew signal tristate
rlabel metal2 s 18786 0 18842 800 6 HI[349]
port 276 nsew signal tristate
rlabel metal2 s 43810 0 43866 800 6 HI[34]
port 277 nsew signal tristate
rlabel metal2 s 5906 3800 5962 4600 6 HI[350]
port 278 nsew signal tristate
rlabel metal2 s 34426 0 34482 800 6 HI[351]
port 279 nsew signal tristate
rlabel metal2 s 48042 3800 48098 4600 6 HI[352]
port 280 nsew signal tristate
rlabel metal2 s 16578 3800 16634 4600 6 HI[353]
port 281 nsew signal tristate
rlabel metal2 s 44914 3800 44970 4600 6 HI[354]
port 282 nsew signal tristate
rlabel metal2 s 6458 3800 6514 4600 6 HI[355]
port 283 nsew signal tristate
rlabel metal2 s 50434 3800 50490 4600 6 HI[356]
port 284 nsew signal tristate
rlabel metal2 s 57242 0 57298 800 6 HI[357]
port 285 nsew signal tristate
rlabel metal2 s 35346 3800 35402 4600 6 HI[358]
port 286 nsew signal tristate
rlabel metal2 s 43626 3800 43682 4600 6 HI[359]
port 287 nsew signal tristate
rlabel metal2 s 54114 3800 54170 4600 6 HI[35]
port 288 nsew signal tristate
rlabel metal2 s 49330 0 49386 800 6 HI[360]
port 289 nsew signal tristate
rlabel metal3 s 59200 1640 60000 1760 6 HI[361]
port 290 nsew signal tristate
rlabel metal2 s 8482 0 8538 800 6 HI[362]
port 291 nsew signal tristate
rlabel metal3 s 59200 1096 60000 1216 6 HI[363]
port 292 nsew signal tristate
rlabel metal2 s 29274 3800 29330 4600 6 HI[364]
port 293 nsew signal tristate
rlabel metal2 s 28354 0 28410 800 6 HI[365]
port 294 nsew signal tristate
rlabel metal2 s 27986 3800 28042 4600 6 HI[366]
port 295 nsew signal tristate
rlabel metal2 s 46938 0 46994 800 6 HI[367]
port 296 nsew signal tristate
rlabel metal2 s 55218 0 55274 800 6 HI[368]
port 297 nsew signal tristate
rlabel metal2 s 51354 0 51410 800 6 HI[369]
port 298 nsew signal tristate
rlabel metal2 s 24306 0 24362 800 6 HI[36]
port 299 nsew signal tristate
rlabel metal2 s 49882 3800 49938 4600 6 HI[370]
port 300 nsew signal tristate
rlabel metal3 s 0 1096 800 1216 6 HI[371]
port 301 nsew signal tristate
rlabel metal2 s 21362 3800 21418 4600 6 HI[372]
port 302 nsew signal tristate
rlabel metal2 s 19338 0 19394 800 6 HI[373]
port 303 nsew signal tristate
rlabel metal2 s 29458 3800 29514 4600 6 HI[374]
port 304 nsew signal tristate
rlabel metal2 s 26514 3800 26570 4600 6 HI[375]
port 305 nsew signal tristate
rlabel metal2 s 53930 3800 53986 4600 6 HI[376]
port 306 nsew signal tristate
rlabel metal2 s 9586 3800 9642 4600 6 HI[377]
port 307 nsew signal tristate
rlabel metal2 s 15842 0 15898 800 6 HI[378]
port 308 nsew signal tristate
rlabel metal2 s 14554 0 14610 800 6 HI[379]
port 309 nsew signal tristate
rlabel metal2 s 16762 3800 16818 4600 6 HI[37]
port 310 nsew signal tristate
rlabel metal2 s 38474 3800 38530 4600 6 HI[380]
port 311 nsew signal tristate
rlabel metal2 s 570 3800 626 4600 6 HI[381]
port 312 nsew signal tristate
rlabel metal2 s 24122 0 24178 800 6 HI[382]
port 313 nsew signal tristate
rlabel metal2 s 6642 3800 6698 4600 6 HI[383]
port 314 nsew signal tristate
rlabel metal2 s 50618 0 50674 800 6 HI[384]
port 315 nsew signal tristate
rlabel metal2 s 30010 3800 30066 4600 6 HI[385]
port 316 nsew signal tristate
rlabel metal2 s 19890 0 19946 800 6 HI[386]
port 317 nsew signal tristate
rlabel metal2 s 45650 3800 45706 4600 6 HI[387]
port 318 nsew signal tristate
rlabel metal2 s 5170 0 5226 800 6 HI[388]
port 319 nsew signal tristate
rlabel metal2 s 31850 3800 31906 4600 6 HI[389]
port 320 nsew signal tristate
rlabel metal2 s 23202 3800 23258 4600 6 HI[38]
port 321 nsew signal tristate
rlabel metal2 s 57794 0 57850 800 6 HI[390]
port 322 nsew signal tristate
rlabel metal2 s 21730 0 21786 800 6 HI[391]
port 323 nsew signal tristate
rlabel metal2 s 26514 0 26570 800 6 HI[392]
port 324 nsew signal tristate
rlabel metal2 s 47490 3800 47546 4600 6 HI[393]
port 325 nsew signal tristate
rlabel metal2 s 44178 0 44234 800 6 HI[394]
port 326 nsew signal tristate
rlabel metal2 s 20994 3800 21050 4600 6 HI[395]
port 327 nsew signal tristate
rlabel metal2 s 57058 3800 57114 4600 6 HI[396]
port 328 nsew signal tristate
rlabel metal2 s 13450 0 13506 800 6 HI[397]
port 329 nsew signal tristate
rlabel metal2 s 28722 3800 28778 4600 6 HI[398]
port 330 nsew signal tristate
rlabel metal2 s 22834 3800 22890 4600 6 HI[399]
port 331 nsew signal tristate
rlabel metal2 s 31482 0 31538 800 6 HI[39]
port 332 nsew signal tristate
rlabel metal2 s 16394 0 16450 800 6 HI[3]
port 333 nsew signal tristate
rlabel metal2 s 32402 0 32458 800 6 HI[400]
port 334 nsew signal tristate
rlabel metal2 s 36634 0 36690 800 6 HI[401]
port 335 nsew signal tristate
rlabel metal2 s 15658 3800 15714 4600 6 HI[402]
port 336 nsew signal tristate
rlabel metal2 s 7562 3800 7618 4600 6 HI[403]
port 337 nsew signal tristate
rlabel metal2 s 56506 3800 56562 4600 6 HI[404]
port 338 nsew signal tristate
rlabel metal2 s 41050 0 41106 800 6 HI[405]
port 339 nsew signal tristate
rlabel metal2 s 48594 0 48650 800 6 HI[406]
port 340 nsew signal tristate
rlabel metal2 s 43994 0 44050 800 6 HI[407]
port 341 nsew signal tristate
rlabel metal2 s 8850 3800 8906 4600 6 HI[408]
port 342 nsew signal tristate
rlabel metal2 s 37554 3800 37610 4600 6 HI[409]
port 343 nsew signal tristate
rlabel metal2 s 20074 0 20130 800 6 HI[40]
port 344 nsew signal tristate
rlabel metal2 s 38474 0 38530 800 6 HI[410]
port 345 nsew signal tristate
rlabel metal2 s 2410 0 2466 800 6 HI[411]
port 346 nsew signal tristate
rlabel metal2 s 55586 0 55642 800 6 HI[412]
port 347 nsew signal tristate
rlabel metal2 s 13266 0 13322 800 6 HI[413]
port 348 nsew signal tristate
rlabel metal2 s 16210 0 16266 800 6 HI[414]
port 349 nsew signal tristate
rlabel metal2 s 29642 0 29698 800 6 HI[415]
port 350 nsew signal tristate
rlabel metal2 s 30378 3800 30434 4600 6 HI[416]
port 351 nsew signal tristate
rlabel metal2 s 35530 0 35586 800 6 HI[417]
port 352 nsew signal tristate
rlabel metal2 s 55770 3800 55826 4600 6 HI[418]
port 353 nsew signal tristate
rlabel metal2 s 30194 0 30250 800 6 HI[419]
port 354 nsew signal tristate
rlabel metal2 s 34242 3800 34298 4600 6 HI[41]
port 355 nsew signal tristate
rlabel metal2 s 33690 0 33746 800 6 HI[420]
port 356 nsew signal tristate
rlabel metal2 s 15106 3800 15162 4600 6 HI[421]
port 357 nsew signal tristate
rlabel metal2 s 11978 3800 12034 4600 6 HI[422]
port 358 nsew signal tristate
rlabel metal2 s 57058 0 57114 800 6 HI[423]
port 359 nsew signal tristate
rlabel metal2 s 35162 0 35218 800 6 HI[424]
port 360 nsew signal tristate
rlabel metal2 s 58162 3800 58218 4600 6 HI[425]
port 361 nsew signal tristate
rlabel metal2 s 9954 3800 10010 4600 6 HI[426]
port 362 nsew signal tristate
rlabel metal2 s 58714 3800 58770 4600 6 HI[427]
port 363 nsew signal tristate
rlabel metal2 s 44730 0 44786 800 6 HI[428]
port 364 nsew signal tristate
rlabel metal3 s 0 3544 800 3664 6 HI[429]
port 365 nsew signal tristate
rlabel metal2 s 1858 0 1914 800 6 HI[42]
port 366 nsew signal tristate
rlabel metal2 s 36082 3800 36138 4600 6 HI[430]
port 367 nsew signal tristate
rlabel metal2 s 34610 3800 34666 4600 6 HI[431]
port 368 nsew signal tristate
rlabel metal2 s 17314 3800 17370 4600 6 HI[432]
port 369 nsew signal tristate
rlabel metal2 s 18050 3800 18106 4600 6 HI[433]
port 370 nsew signal tristate
rlabel metal2 s 48410 3800 48466 4600 6 HI[434]
port 371 nsew signal tristate
rlabel metal2 s 16210 3800 16266 4600 6 HI[435]
port 372 nsew signal tristate
rlabel metal2 s 16946 0 17002 800 6 HI[436]
port 373 nsew signal tristate
rlabel metal2 s 18234 0 18290 800 6 HI[437]
port 374 nsew signal tristate
rlabel metal2 s 55034 3800 55090 4600 6 HI[438]
port 375 nsew signal tristate
rlabel metal3 s 59200 2728 60000 2848 6 HI[439]
port 376 nsew signal tristate
rlabel metal2 s 2042 0 2098 800 6 HI[43]
port 377 nsew signal tristate
rlabel metal2 s 20994 0 21050 800 6 HI[440]
port 378 nsew signal tristate
rlabel metal2 s 46754 3800 46810 4600 6 HI[441]
port 379 nsew signal tristate
rlabel metal2 s 13818 3800 13874 4600 6 HI[442]
port 380 nsew signal tristate
rlabel metal2 s 52090 3800 52146 4600 6 HI[443]
port 381 nsew signal tristate
rlabel metal2 s 14186 3800 14242 4600 6 HI[444]
port 382 nsew signal tristate
rlabel metal2 s 25778 3800 25834 4600 6 HI[445]
port 383 nsew signal tristate
rlabel metal2 s 31850 0 31906 800 6 HI[446]
port 384 nsew signal tristate
rlabel metal2 s 21914 0 21970 800 6 HI[447]
port 385 nsew signal tristate
rlabel metal2 s 10322 0 10378 800 6 HI[448]
port 386 nsew signal tristate
rlabel metal2 s 1490 0 1546 800 6 HI[449]
port 387 nsew signal tristate
rlabel metal2 s 8298 3800 8354 4600 6 HI[44]
port 388 nsew signal tristate
rlabel metal2 s 18418 3800 18474 4600 6 HI[450]
port 389 nsew signal tristate
rlabel metal2 s 55954 0 56010 800 6 HI[451]
port 390 nsew signal tristate
rlabel metal2 s 27802 0 27858 800 6 HI[452]
port 391 nsew signal tristate
rlabel metal2 s 5538 3800 5594 4600 6 HI[453]
port 392 nsew signal tristate
rlabel metal2 s 24490 3800 24546 4600 6 HI[454]
port 393 nsew signal tristate
rlabel metal2 s 30930 0 30986 800 6 HI[455]
port 394 nsew signal tristate
rlabel metal2 s 48962 0 49018 800 6 HI[456]
port 395 nsew signal tristate
rlabel metal2 s 17866 3800 17922 4600 6 HI[457]
port 396 nsew signal tristate
rlabel metal2 s 45650 0 45706 800 6 HI[458]
port 397 nsew signal tristate
rlabel metal2 s 40314 3800 40370 4600 6 HI[45]
port 398 nsew signal tristate
rlabel metal2 s 51722 0 51778 800 6 HI[46]
port 399 nsew signal tristate
rlabel metal2 s 7194 0 7250 800 6 HI[47]
port 400 nsew signal tristate
rlabel metal2 s 51906 0 51962 800 6 HI[48]
port 401 nsew signal tristate
rlabel metal2 s 30746 3800 30802 4600 6 HI[49]
port 402 nsew signal tristate
rlabel metal2 s 39210 0 39266 800 6 HI[4]
port 403 nsew signal tristate
rlabel metal2 s 56138 0 56194 800 6 HI[50]
port 404 nsew signal tristate
rlabel metal2 s 57610 0 57666 800 6 HI[51]
port 405 nsew signal tristate
rlabel metal2 s 48962 3800 49018 4600 6 HI[52]
port 406 nsew signal tristate
rlabel metal2 s 20258 3800 20314 4600 6 HI[53]
port 407 nsew signal tristate
rlabel metal2 s 57426 3800 57482 4600 6 HI[54]
port 408 nsew signal tristate
rlabel metal2 s 59082 0 59138 800 6 HI[55]
port 409 nsew signal tristate
rlabel metal2 s 21178 0 21234 800 6 HI[56]
port 410 nsew signal tristate
rlabel metal2 s 55954 3800 56010 4600 6 HI[57]
port 411 nsew signal tristate
rlabel metal2 s 19338 3800 19394 4600 6 HI[58]
port 412 nsew signal tristate
rlabel metal2 s 52826 0 52882 800 6 HI[59]
port 413 nsew signal tristate
rlabel metal2 s 35162 3800 35218 4600 6 HI[5]
port 414 nsew signal tristate
rlabel metal2 s 50250 3800 50306 4600 6 HI[60]
port 415 nsew signal tristate
rlabel metal2 s 20626 0 20682 800 6 HI[61]
port 416 nsew signal tristate
rlabel metal2 s 13818 0 13874 800 6 HI[62]
port 417 nsew signal tristate
rlabel metal2 s 48042 0 48098 800 6 HI[63]
port 418 nsew signal tristate
rlabel metal2 s 24858 0 24914 800 6 HI[64]
port 419 nsew signal tristate
rlabel metal2 s 50986 0 51042 800 6 HI[65]
port 420 nsew signal tristate
rlabel metal2 s 25226 0 25282 800 6 HI[66]
port 421 nsew signal tristate
rlabel metal2 s 33138 0 33194 800 6 HI[67]
port 422 nsew signal tristate
rlabel metal2 s 754 0 810 800 6 HI[68]
port 423 nsew signal tristate
rlabel metal2 s 41418 0 41474 800 6 HI[69]
port 424 nsew signal tristate
rlabel metal2 s 46570 0 46626 800 6 HI[6]
port 425 nsew signal tristate
rlabel metal2 s 3514 3800 3570 4600 6 HI[70]
port 426 nsew signal tristate
rlabel metal3 s 0 2728 800 2848 6 HI[71]
port 427 nsew signal tristate
rlabel metal2 s 4066 3800 4122 4600 6 HI[72]
port 428 nsew signal tristate
rlabel metal2 s 13634 3800 13690 4600 6 HI[73]
port 429 nsew signal tristate
rlabel metal2 s 21362 0 21418 800 6 HI[74]
port 430 nsew signal tristate
rlabel metal2 s 49698 3800 49754 4600 6 HI[75]
port 431 nsew signal tristate
rlabel metal2 s 44546 3800 44602 4600 6 HI[76]
port 432 nsew signal tristate
rlabel metal2 s 33506 3800 33562 4600 6 HI[77]
port 433 nsew signal tristate
rlabel metal2 s 49146 3800 49202 4600 6 HI[78]
port 434 nsew signal tristate
rlabel metal2 s 46570 3800 46626 4600 6 HI[79]
port 435 nsew signal tristate
rlabel metal2 s 49514 0 49570 800 6 HI[7]
port 436 nsew signal tristate
rlabel metal2 s 32218 3800 32274 4600 6 HI[80]
port 437 nsew signal tristate
rlabel metal2 s 51354 3800 51410 4600 6 HI[81]
port 438 nsew signal tristate
rlabel metal2 s 57978 0 58034 800 6 HI[82]
port 439 nsew signal tristate
rlabel metal2 s 17498 3800 17554 4600 6 HI[83]
port 440 nsew signal tristate
rlabel metal2 s 20810 3800 20866 4600 6 HI[84]
port 441 nsew signal tristate
rlabel metal2 s 10138 3800 10194 4600 6 HI[85]
port 442 nsew signal tristate
rlabel metal2 s 31114 3800 31170 4600 6 HI[86]
port 443 nsew signal tristate
rlabel metal2 s 22466 0 22522 800 6 HI[87]
port 444 nsew signal tristate
rlabel metal2 s 53194 3800 53250 4600 6 HI[88]
port 445 nsew signal tristate
rlabel metal2 s 1858 3800 1914 4600 6 HI[89]
port 446 nsew signal tristate
rlabel metal2 s 37922 3800 37978 4600 6 HI[8]
port 447 nsew signal tristate
rlabel metal2 s 1122 3800 1178 4600 6 HI[90]
port 448 nsew signal tristate
rlabel metal2 s 26882 3800 26938 4600 6 HI[91]
port 449 nsew signal tristate
rlabel metal2 s 3146 3800 3202 4600 6 HI[92]
port 450 nsew signal tristate
rlabel metal2 s 29090 0 29146 800 6 HI[93]
port 451 nsew signal tristate
rlabel metal2 s 46018 3800 46074 4600 6 HI[94]
port 452 nsew signal tristate
rlabel metal2 s 2778 3800 2834 4600 6 HI[95]
port 453 nsew signal tristate
rlabel metal2 s 17682 0 17738 800 6 HI[96]
port 454 nsew signal tristate
rlabel metal2 s 15474 3800 15530 4600 6 HI[97]
port 455 nsew signal tristate
rlabel metal2 s 25962 0 26018 800 6 HI[98]
port 456 nsew signal tristate
rlabel metal3 s 59200 824 60000 944 6 HI[99]
port 457 nsew signal tristate
rlabel metal2 s 36266 0 36322 800 6 HI[9]
port 458 nsew signal tristate
rlabel metal2 s 51350 1040 51410 3312 6 vccd1
port 459 nsew power bidirectional
rlabel metal2 s 35350 1040 35410 3312 6 vccd1
port 460 nsew power bidirectional
rlabel metal2 s 19350 1040 19410 3312 6 vccd1
port 461 nsew power bidirectional
rlabel metal2 s 3350 1040 3410 3312 6 vccd1
port 462 nsew power bidirectional
rlabel metal3 s 1380 1210 58604 1270 6 vccd1
port 463 nsew power bidirectional
rlabel metal2 s 43350 1040 43410 3312 6 vssd1
port 464 nsew ground bidirectional
rlabel metal2 s 27350 1040 27410 3312 6 vssd1
port 465 nsew ground bidirectional
rlabel metal2 s 11350 1040 11410 3312 6 vssd1
port 466 nsew ground bidirectional
rlabel metal3 s 1380 2290 58604 2350 6 vssd1
port 467 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 4600
<< end >>
