magic
tech sky130A
magscale 1 2
timestamp 1661898952
<< nwell >>
rect 530 550 1000 890
rect 590 -980 930 550
<< pmoslvt >>
rect 720 320 820 520
rect 720 0 820 200
rect 730 -870 800 -270
<< nmoslvt >>
rect 770 -1260 800 -1060
rect 710 -2220 740 -1420
rect 820 -2220 850 -1420
rect 730 -2660 830 -2460
<< ndiff >>
rect 700 -1080 770 -1060
rect 700 -1240 710 -1080
rect 750 -1240 770 -1080
rect 700 -1260 770 -1240
rect 800 -1080 870 -1060
rect 800 -1240 820 -1080
rect 860 -1240 870 -1080
rect 800 -1260 870 -1240
rect 640 -1420 690 -1380
rect 640 -1440 710 -1420
rect 640 -2200 650 -1440
rect 690 -2200 710 -1440
rect 640 -2220 710 -2200
rect 740 -1440 820 -1420
rect 740 -2200 760 -1440
rect 800 -2200 820 -1440
rect 740 -2220 820 -2200
rect 850 -1440 920 -1420
rect 850 -2190 870 -1440
rect 910 -2190 920 -1440
rect 850 -2220 920 -2190
rect 730 -2400 830 -2390
rect 730 -2440 750 -2400
rect 810 -2440 830 -2400
rect 730 -2460 830 -2440
rect 730 -2710 830 -2660
rect 730 -2750 750 -2710
rect 810 -2750 830 -2710
rect 730 -2760 830 -2750
<< pdiff >>
rect 640 500 720 520
rect 640 340 660 500
rect 700 340 720 500
rect 640 320 720 340
rect 820 500 890 520
rect 820 340 840 500
rect 880 340 890 500
rect 820 320 890 340
rect 650 180 720 200
rect 650 20 660 180
rect 700 20 720 180
rect 650 0 720 20
rect 820 180 890 200
rect 820 20 840 180
rect 880 20 890 180
rect 820 0 890 20
rect 660 -290 730 -270
rect 660 -850 670 -290
rect 710 -850 730 -290
rect 660 -870 730 -850
rect 800 -290 870 -270
rect 800 -850 820 -290
rect 860 -850 870 -290
rect 800 -870 870 -850
<< ndiffc >>
rect 710 -1240 750 -1080
rect 820 -1240 860 -1080
rect 650 -2200 690 -1440
rect 760 -2200 800 -1440
rect 870 -2190 910 -1440
rect 750 -2440 810 -2400
rect 750 -2750 810 -2710
<< pdiffc >>
rect 660 340 700 500
rect 840 340 880 500
rect 660 20 700 180
rect 840 20 880 180
rect 670 -850 710 -290
rect 820 -850 860 -290
<< psubdiff >>
rect 590 -2840 930 -2820
rect 590 -2890 660 -2840
rect 900 -2890 930 -2840
rect 590 -2900 930 -2890
<< nsubdiff >>
rect 640 750 720 780
rect 590 610 620 750
rect 870 610 930 750
rect 640 580 720 610
<< psubdiffcont >>
rect 660 -2890 900 -2840
<< nsubdiffcont >>
rect 620 610 870 750
<< poly >>
rect 720 520 820 550
rect 720 200 820 320
rect 720 -30 820 0
rect 750 -40 820 -30
rect 750 -53 830 -40
rect 750 -87 783 -53
rect 817 -87 830 -53
rect 750 -120 830 -87
rect 730 -180 810 -170
rect 730 -220 750 -180
rect 790 -220 810 -180
rect 730 -230 810 -220
rect 730 -270 800 -230
rect 730 -1000 800 -870
rect 770 -1060 800 -1000
rect 770 -1290 800 -1260
rect 710 -1420 740 -1390
rect 820 -1420 850 -1390
rect 710 -2280 740 -2220
rect 630 -2298 740 -2280
rect 630 -2332 653 -2298
rect 687 -2332 740 -2298
rect 630 -2350 740 -2332
rect 820 -2280 850 -2220
rect 820 -2298 920 -2280
rect 820 -2332 873 -2298
rect 907 -2332 920 -2298
rect 820 -2350 920 -2332
rect 700 -2600 730 -2460
rect 630 -2610 730 -2600
rect 630 -2650 650 -2610
rect 690 -2650 730 -2610
rect 630 -2660 730 -2650
rect 830 -2660 860 -2460
<< polycont >>
rect 783 -87 817 -53
rect 750 -220 790 -180
rect 653 -2332 687 -2298
rect 873 -2332 907 -2298
rect 650 -2650 690 -2610
<< locali >>
rect 640 750 720 780
rect 590 730 620 750
rect 870 730 930 750
rect 590 630 600 730
rect 890 630 930 730
rect 590 610 620 630
rect 870 610 930 630
rect 640 580 720 610
rect 650 500 700 580
rect 650 340 660 500
rect 650 320 700 340
rect 840 500 880 520
rect 660 180 700 320
rect 660 -270 700 20
rect 840 180 890 200
rect 880 20 890 180
rect 840 -50 890 20
rect 750 -52 890 -50
rect 784 -53 890 -52
rect 750 -87 783 -86
rect 817 -87 890 -53
rect 750 -90 890 -87
rect 750 -180 790 -160
rect 740 -220 750 -180
rect 790 -183 810 -180
rect 797 -217 810 -183
rect 790 -220 810 -217
rect 850 -220 890 -90
rect 750 -240 790 -220
rect 660 -290 710 -270
rect 660 -850 670 -290
rect 660 -870 710 -850
rect 820 -290 870 -270
rect 860 -850 870 -290
rect 820 -970 860 -850
rect 810 -1010 860 -970
rect 700 -1080 760 -1060
rect 700 -1240 710 -1080
rect 750 -1090 760 -1080
rect 700 -1260 760 -1240
rect 820 -1080 860 -1010
rect 820 -1260 860 -1240
rect 630 -1440 700 -1380
rect 630 -2200 640 -1440
rect 690 -2200 700 -1440
rect 630 -2220 700 -2200
rect 760 -1440 800 -1390
rect 653 -2298 687 -2282
rect 653 -2348 687 -2332
rect 760 -2390 800 -2200
rect 860 -1440 920 -1420
rect 860 -1460 870 -1440
rect 910 -2190 920 -1440
rect 900 -2200 920 -2190
rect 860 -2220 920 -2200
rect 873 -2298 907 -2282
rect 873 -2348 907 -2332
rect 730 -2400 830 -2390
rect 730 -2440 750 -2400
rect 810 -2440 830 -2400
rect 630 -2600 710 -2590
rect 630 -2660 640 -2600
rect 700 -2660 710 -2600
rect 630 -2670 710 -2660
rect 730 -2710 830 -2700
rect 730 -2750 750 -2710
rect 810 -2750 830 -2710
rect 730 -2820 830 -2750
rect 590 -2840 930 -2820
rect 590 -2890 660 -2840
rect 900 -2890 930 -2840
rect 590 -2900 930 -2890
<< viali >>
rect 600 630 620 730
rect 620 630 870 730
rect 870 630 890 730
rect 840 340 880 470
rect 840 320 880 340
rect 750 -53 784 -52
rect 750 -86 783 -53
rect 783 -86 784 -53
rect 763 -217 790 -183
rect 790 -217 797 -183
rect 770 -1010 810 -970
rect 720 -1240 750 -1090
rect 750 -1240 760 -1090
rect 640 -2200 650 -1440
rect 650 -2200 680 -1440
rect 653 -2332 687 -2298
rect 860 -2190 870 -1460
rect 870 -2190 900 -1460
rect 860 -2200 900 -2190
rect 873 -2332 907 -2298
rect 640 -2610 700 -2600
rect 640 -2650 650 -2610
rect 650 -2650 690 -2610
rect 690 -2650 700 -2610
rect 640 -2660 700 -2650
rect 660 -2890 900 -2840
<< metal1 >>
rect 590 730 930 780
rect 590 630 600 730
rect 890 630 930 730
rect 590 580 930 630
rect 830 470 890 490
rect 830 320 840 470
rect 880 320 890 470
rect 830 290 890 320
rect 630 -52 670 -50
rect 744 -52 790 -40
rect 630 -85 750 -52
rect 630 -1380 670 -85
rect 744 -86 750 -85
rect 784 -86 790 -52
rect 744 -98 790 -86
rect 830 -170 860 290
rect 740 -183 860 -170
rect 740 -217 763 -183
rect 797 -217 860 -183
rect 740 -230 860 -217
rect 750 -250 790 -230
rect 820 -235 860 -230
rect 820 -270 905 -235
rect 764 -964 816 -958
rect 764 -1022 816 -1016
rect 710 -1090 770 -1060
rect 710 -1240 720 -1090
rect 760 -1240 770 -1090
rect 710 -1260 780 -1240
rect 740 -1298 780 -1260
rect 734 -1304 786 -1298
rect 875 -1320 905 -270
rect 734 -1362 786 -1356
rect 630 -1440 700 -1380
rect 630 -2200 640 -1440
rect 680 -2200 700 -1440
rect 630 -2220 700 -2200
rect 850 -1460 910 -1320
rect 850 -2200 860 -1460
rect 900 -2200 910 -1460
rect 850 -2220 910 -2200
rect 644 -2289 696 -2283
rect 644 -2347 696 -2341
rect 864 -2289 916 -2283
rect 864 -2347 916 -2341
rect 634 -2590 706 -2588
rect 630 -2600 790 -2590
rect 630 -2660 640 -2600
rect 700 -2660 720 -2600
rect 780 -2660 790 -2600
rect 630 -2670 790 -2660
rect 634 -2672 706 -2670
rect 590 -2830 930 -2790
rect 590 -2840 680 -2830
rect 880 -2840 930 -2830
rect 590 -2890 660 -2840
rect 900 -2890 930 -2840
rect 590 -2990 930 -2890
<< via1 >>
rect 764 -970 816 -964
rect 764 -1010 770 -970
rect 770 -1010 810 -970
rect 810 -1010 816 -970
rect 764 -1016 816 -1010
rect 734 -1356 786 -1304
rect 644 -2298 696 -2289
rect 644 -2332 653 -2298
rect 653 -2332 687 -2298
rect 687 -2332 696 -2298
rect 644 -2341 696 -2332
rect 864 -2298 916 -2289
rect 864 -2332 873 -2298
rect 873 -2332 907 -2298
rect 907 -2332 916 -2298
rect 864 -2341 916 -2332
rect 720 -2660 780 -2600
rect 680 -2840 880 -2830
rect 680 -2890 880 -2840
<< metal2 >>
rect 750 -960 830 -950
rect 750 -1020 760 -960
rect 820 -1020 830 -960
rect 750 -1030 830 -1020
rect 728 -1356 734 -1304
rect 786 -1310 792 -1304
rect 786 -1356 800 -1310
rect 630 -2340 640 -2280
rect 700 -2340 710 -2280
rect 630 -2341 644 -2340
rect 696 -2341 710 -2340
rect 630 -2350 710 -2341
rect 760 -2520 800 -1356
rect 873 -2289 907 977
rect 858 -2341 864 -2289
rect 916 -2341 922 -2289
rect 640 -2560 800 -2520
rect 640 -2820 680 -2560
rect 710 -2600 800 -2590
rect 710 -2660 720 -2600
rect 780 -2660 800 -2600
rect 710 -2670 800 -2660
rect 640 -2830 900 -2820
rect 640 -2890 680 -2830
rect 880 -2890 900 -2830
rect 640 -2900 900 -2890
<< via2 >>
rect 760 -964 820 -960
rect 760 -1016 764 -964
rect 764 -1016 816 -964
rect 816 -1016 820 -964
rect 760 -1020 820 -1016
rect 640 -2289 700 -2280
rect 640 -2340 644 -2289
rect 644 -2340 696 -2289
rect 696 -2340 700 -2289
rect 720 -2660 780 -2600
<< metal3 >>
rect 740 -955 840 -940
rect 740 -1025 755 -955
rect 825 -1025 840 -955
rect 740 -1040 840 -1025
rect 630 -2280 710 -2270
rect 630 -2340 640 -2280
rect 700 -2340 970 -2280
rect 630 -2350 970 -2340
rect 715 -2600 785 -2595
rect 590 -2660 720 -2600
rect 780 -2660 930 -2600
rect 715 -2665 785 -2660
<< via3 >>
rect 755 -960 825 -955
rect 755 -1020 760 -960
rect 760 -1020 820 -960
rect 820 -1020 825 -960
rect 755 -1025 825 -1020
<< metal4 >>
rect 750 -955 830 -950
rect 750 -1025 755 -955
rect 825 -1025 830 -955
rect 750 -1030 830 -1025
rect 760 -3100 820 -1030
<< labels >>
rlabel metal2 890 940 890 940 1 V_IN
port 1 n
rlabel metal1 600 600 600 600 1 VDD
port 2 n
rlabel metal1 660 -2940 660 -2940 1 GND
port 3 n
rlabel metal3 600 -2630 600 -2630 1 SA_IREF
port 5 n
rlabel metal4 790 -3000 790 -3000 1 OUT
port 6 n
rlabel metal1 720 -70 720 -70 1 GN
rlabel metal1 850 270 850 270 1 net1
rlabel locali 740 -2420 740 -2420 1 net2
rlabel metal3 950 -2310 950 -2310 1 REF
port 7 n
<< end >>
