* SPICE3 file created from 8bit_dram.ext - technology: sky130A

.subckt dram_cell WWL WBL RWL RBL VSUBS
X0 RWL storage RBL VSUBS sky130_fd_pr__nfet_01v8 ad=3e+11p pd=2.6e+06u as=3.5e+11p ps=2.7e+06u w=1e+06u l=150000u
X1 storage WWL WBL VSUBS sky130_fd_pr__nfet_01v8 ad=3.5e+11p pd=2.7e+06u as=3e+11p ps=2.6e+06u w=1e+06u l=150000u
.ends

.subckt dram_array READ_BOT READ_TOP WWL WRITE dram_cell_0/WBL dram_cell_1/RWL VSUBS
Xdram_cell_0 WWL dram_cell_0/WBL dram_cell_1/RWL READ_TOP VSUBS dram_cell
Xdram_cell_1 WWL WRITE dram_cell_1/RWL READ_BOT VSUBS dram_cell
.ends

.subckt x4bit_dram dram_array_1/READ_TOP dram_array_1/READ_BOT dram_array_0/WRITE
+ dram_array_1/dram_cell_0/WBL dram_array_1/WRITE dram_array_0/dram_cell_0/WBL dram_array_1/dram_cell_1/RWL
+ dram_array_0/READ_TOP dram_array_0/READ_BOT dram_array_1/WWL VSUBS
Xdram_array_0 dram_array_0/READ_BOT dram_array_0/READ_TOP dram_array_1/WWL dram_array_0/WRITE
+ dram_array_0/dram_cell_0/WBL dram_array_1/dram_cell_1/RWL VSUBS dram_array
Xdram_array_1 dram_array_1/READ_BOT dram_array_1/READ_TOP dram_array_1/WWL dram_array_1/WRITE
+ dram_array_1/dram_cell_0/WBL dram_array_1/dram_cell_1/RWL VSUBS dram_array
.ends

.subckt x8bit_dram READ WRITE INx0x OUTx0x OUTX4x INx1x OUTx1x OUTx5x INx2x OUTx2x
+ OUTx6x INx3x OUTx7x OUTx3x INx4x INx5x INx6x INx7x
X4bit_dram_1 OUTx3x OUTx7x INx6x INx3x INx7x INx2x READ OUTx2x OUTx6x WRITE VSUBS
+ x4bit_dram
X4bit_dram_0 OUTx1x OUTx5x INx4x INx1x INx5x INx0x READ OUTx0x OUTX4x WRITE VSUBS
+ x4bit_dram
.ends

