magic
tech sky130B
magscale 1 2
timestamp 1607714484
<< pwell >>
rect -1947 -1519 1947 1519
<< nmos >>
rect -1751 109 -1631 1309
rect -1573 109 -1453 1309
rect -1395 109 -1275 1309
rect -1217 109 -1097 1309
rect -1039 109 -919 1309
rect -861 109 -741 1309
rect -683 109 -563 1309
rect -505 109 -385 1309
rect -327 109 -207 1309
rect -149 109 -29 1309
rect 29 109 149 1309
rect 207 109 327 1309
rect 385 109 505 1309
rect 563 109 683 1309
rect 741 109 861 1309
rect 919 109 1039 1309
rect 1097 109 1217 1309
rect 1275 109 1395 1309
rect 1453 109 1573 1309
rect 1631 109 1751 1309
rect -1751 -1309 -1631 -109
rect -1573 -1309 -1453 -109
rect -1395 -1309 -1275 -109
rect -1217 -1309 -1097 -109
rect -1039 -1309 -919 -109
rect -861 -1309 -741 -109
rect -683 -1309 -563 -109
rect -505 -1309 -385 -109
rect -327 -1309 -207 -109
rect -149 -1309 -29 -109
rect 29 -1309 149 -109
rect 207 -1309 327 -109
rect 385 -1309 505 -109
rect 563 -1309 683 -109
rect 741 -1309 861 -109
rect 919 -1309 1039 -109
rect 1097 -1309 1217 -109
rect 1275 -1309 1395 -109
rect 1453 -1309 1573 -109
rect 1631 -1309 1751 -109
<< ndiff >>
rect -1809 1297 -1751 1309
rect -1809 121 -1797 1297
rect -1763 121 -1751 1297
rect -1809 109 -1751 121
rect -1631 1297 -1573 1309
rect -1631 121 -1619 1297
rect -1585 121 -1573 1297
rect -1631 109 -1573 121
rect -1453 1297 -1395 1309
rect -1453 121 -1441 1297
rect -1407 121 -1395 1297
rect -1453 109 -1395 121
rect -1275 1297 -1217 1309
rect -1275 121 -1263 1297
rect -1229 121 -1217 1297
rect -1275 109 -1217 121
rect -1097 1297 -1039 1309
rect -1097 121 -1085 1297
rect -1051 121 -1039 1297
rect -1097 109 -1039 121
rect -919 1297 -861 1309
rect -919 121 -907 1297
rect -873 121 -861 1297
rect -919 109 -861 121
rect -741 1297 -683 1309
rect -741 121 -729 1297
rect -695 121 -683 1297
rect -741 109 -683 121
rect -563 1297 -505 1309
rect -563 121 -551 1297
rect -517 121 -505 1297
rect -563 109 -505 121
rect -385 1297 -327 1309
rect -385 121 -373 1297
rect -339 121 -327 1297
rect -385 109 -327 121
rect -207 1297 -149 1309
rect -207 121 -195 1297
rect -161 121 -149 1297
rect -207 109 -149 121
rect -29 1297 29 1309
rect -29 121 -17 1297
rect 17 121 29 1297
rect -29 109 29 121
rect 149 1297 207 1309
rect 149 121 161 1297
rect 195 121 207 1297
rect 149 109 207 121
rect 327 1297 385 1309
rect 327 121 339 1297
rect 373 121 385 1297
rect 327 109 385 121
rect 505 1297 563 1309
rect 505 121 517 1297
rect 551 121 563 1297
rect 505 109 563 121
rect 683 1297 741 1309
rect 683 121 695 1297
rect 729 121 741 1297
rect 683 109 741 121
rect 861 1297 919 1309
rect 861 121 873 1297
rect 907 121 919 1297
rect 861 109 919 121
rect 1039 1297 1097 1309
rect 1039 121 1051 1297
rect 1085 121 1097 1297
rect 1039 109 1097 121
rect 1217 1297 1275 1309
rect 1217 121 1229 1297
rect 1263 121 1275 1297
rect 1217 109 1275 121
rect 1395 1297 1453 1309
rect 1395 121 1407 1297
rect 1441 121 1453 1297
rect 1395 109 1453 121
rect 1573 1297 1631 1309
rect 1573 121 1585 1297
rect 1619 121 1631 1297
rect 1573 109 1631 121
rect 1751 1297 1809 1309
rect 1751 121 1763 1297
rect 1797 121 1809 1297
rect 1751 109 1809 121
rect -1809 -121 -1751 -109
rect -1809 -1297 -1797 -121
rect -1763 -1297 -1751 -121
rect -1809 -1309 -1751 -1297
rect -1631 -121 -1573 -109
rect -1631 -1297 -1619 -121
rect -1585 -1297 -1573 -121
rect -1631 -1309 -1573 -1297
rect -1453 -121 -1395 -109
rect -1453 -1297 -1441 -121
rect -1407 -1297 -1395 -121
rect -1453 -1309 -1395 -1297
rect -1275 -121 -1217 -109
rect -1275 -1297 -1263 -121
rect -1229 -1297 -1217 -121
rect -1275 -1309 -1217 -1297
rect -1097 -121 -1039 -109
rect -1097 -1297 -1085 -121
rect -1051 -1297 -1039 -121
rect -1097 -1309 -1039 -1297
rect -919 -121 -861 -109
rect -919 -1297 -907 -121
rect -873 -1297 -861 -121
rect -919 -1309 -861 -1297
rect -741 -121 -683 -109
rect -741 -1297 -729 -121
rect -695 -1297 -683 -121
rect -741 -1309 -683 -1297
rect -563 -121 -505 -109
rect -563 -1297 -551 -121
rect -517 -1297 -505 -121
rect -563 -1309 -505 -1297
rect -385 -121 -327 -109
rect -385 -1297 -373 -121
rect -339 -1297 -327 -121
rect -385 -1309 -327 -1297
rect -207 -121 -149 -109
rect -207 -1297 -195 -121
rect -161 -1297 -149 -121
rect -207 -1309 -149 -1297
rect -29 -121 29 -109
rect -29 -1297 -17 -121
rect 17 -1297 29 -121
rect -29 -1309 29 -1297
rect 149 -121 207 -109
rect 149 -1297 161 -121
rect 195 -1297 207 -121
rect 149 -1309 207 -1297
rect 327 -121 385 -109
rect 327 -1297 339 -121
rect 373 -1297 385 -121
rect 327 -1309 385 -1297
rect 505 -121 563 -109
rect 505 -1297 517 -121
rect 551 -1297 563 -121
rect 505 -1309 563 -1297
rect 683 -121 741 -109
rect 683 -1297 695 -121
rect 729 -1297 741 -121
rect 683 -1309 741 -1297
rect 861 -121 919 -109
rect 861 -1297 873 -121
rect 907 -1297 919 -121
rect 861 -1309 919 -1297
rect 1039 -121 1097 -109
rect 1039 -1297 1051 -121
rect 1085 -1297 1097 -121
rect 1039 -1309 1097 -1297
rect 1217 -121 1275 -109
rect 1217 -1297 1229 -121
rect 1263 -1297 1275 -121
rect 1217 -1309 1275 -1297
rect 1395 -121 1453 -109
rect 1395 -1297 1407 -121
rect 1441 -1297 1453 -121
rect 1395 -1309 1453 -1297
rect 1573 -121 1631 -109
rect 1573 -1297 1585 -121
rect 1619 -1297 1631 -121
rect 1573 -1309 1631 -1297
rect 1751 -121 1809 -109
rect 1751 -1297 1763 -121
rect 1797 -1297 1809 -121
rect 1751 -1309 1809 -1297
<< ndiffc >>
rect -1797 121 -1763 1297
rect -1619 121 -1585 1297
rect -1441 121 -1407 1297
rect -1263 121 -1229 1297
rect -1085 121 -1051 1297
rect -907 121 -873 1297
rect -729 121 -695 1297
rect -551 121 -517 1297
rect -373 121 -339 1297
rect -195 121 -161 1297
rect -17 121 17 1297
rect 161 121 195 1297
rect 339 121 373 1297
rect 517 121 551 1297
rect 695 121 729 1297
rect 873 121 907 1297
rect 1051 121 1085 1297
rect 1229 121 1263 1297
rect 1407 121 1441 1297
rect 1585 121 1619 1297
rect 1763 121 1797 1297
rect -1797 -1297 -1763 -121
rect -1619 -1297 -1585 -121
rect -1441 -1297 -1407 -121
rect -1263 -1297 -1229 -121
rect -1085 -1297 -1051 -121
rect -907 -1297 -873 -121
rect -729 -1297 -695 -121
rect -551 -1297 -517 -121
rect -373 -1297 -339 -121
rect -195 -1297 -161 -121
rect -17 -1297 17 -121
rect 161 -1297 195 -121
rect 339 -1297 373 -121
rect 517 -1297 551 -121
rect 695 -1297 729 -121
rect 873 -1297 907 -121
rect 1051 -1297 1085 -121
rect 1229 -1297 1263 -121
rect 1407 -1297 1441 -121
rect 1585 -1297 1619 -121
rect 1763 -1297 1797 -121
<< psubdiff >>
rect -1911 1449 -1815 1483
rect 1815 1449 1911 1483
rect -1911 1387 -1877 1449
rect 1877 1387 1911 1449
rect -1911 -1449 -1877 -1387
rect 1877 -1449 1911 -1387
rect -1911 -1483 -1815 -1449
rect 1815 -1483 1911 -1449
<< psubdiffcont >>
rect -1815 1449 1815 1483
rect -1911 -1387 -1877 1387
rect 1877 -1387 1911 1387
rect -1815 -1483 1815 -1449
<< poly >>
rect -1751 1381 -1631 1397
rect -1751 1347 -1735 1381
rect -1647 1347 -1631 1381
rect -1751 1309 -1631 1347
rect -1573 1381 -1453 1397
rect -1573 1347 -1557 1381
rect -1469 1347 -1453 1381
rect -1573 1309 -1453 1347
rect -1395 1381 -1275 1397
rect -1395 1347 -1379 1381
rect -1291 1347 -1275 1381
rect -1395 1309 -1275 1347
rect -1217 1381 -1097 1397
rect -1217 1347 -1201 1381
rect -1113 1347 -1097 1381
rect -1217 1309 -1097 1347
rect -1039 1381 -919 1397
rect -1039 1347 -1023 1381
rect -935 1347 -919 1381
rect -1039 1309 -919 1347
rect -861 1381 -741 1397
rect -861 1347 -845 1381
rect -757 1347 -741 1381
rect -861 1309 -741 1347
rect -683 1381 -563 1397
rect -683 1347 -667 1381
rect -579 1347 -563 1381
rect -683 1309 -563 1347
rect -505 1381 -385 1397
rect -505 1347 -489 1381
rect -401 1347 -385 1381
rect -505 1309 -385 1347
rect -327 1381 -207 1397
rect -327 1347 -311 1381
rect -223 1347 -207 1381
rect -327 1309 -207 1347
rect -149 1381 -29 1397
rect -149 1347 -133 1381
rect -45 1347 -29 1381
rect -149 1309 -29 1347
rect 29 1381 149 1397
rect 29 1347 45 1381
rect 133 1347 149 1381
rect 29 1309 149 1347
rect 207 1381 327 1397
rect 207 1347 223 1381
rect 311 1347 327 1381
rect 207 1309 327 1347
rect 385 1381 505 1397
rect 385 1347 401 1381
rect 489 1347 505 1381
rect 385 1309 505 1347
rect 563 1381 683 1397
rect 563 1347 579 1381
rect 667 1347 683 1381
rect 563 1309 683 1347
rect 741 1381 861 1397
rect 741 1347 757 1381
rect 845 1347 861 1381
rect 741 1309 861 1347
rect 919 1381 1039 1397
rect 919 1347 935 1381
rect 1023 1347 1039 1381
rect 919 1309 1039 1347
rect 1097 1381 1217 1397
rect 1097 1347 1113 1381
rect 1201 1347 1217 1381
rect 1097 1309 1217 1347
rect 1275 1381 1395 1397
rect 1275 1347 1291 1381
rect 1379 1347 1395 1381
rect 1275 1309 1395 1347
rect 1453 1381 1573 1397
rect 1453 1347 1469 1381
rect 1557 1347 1573 1381
rect 1453 1309 1573 1347
rect 1631 1381 1751 1397
rect 1631 1347 1647 1381
rect 1735 1347 1751 1381
rect 1631 1309 1751 1347
rect -1751 71 -1631 109
rect -1751 37 -1735 71
rect -1647 37 -1631 71
rect -1751 21 -1631 37
rect -1573 71 -1453 109
rect -1573 37 -1557 71
rect -1469 37 -1453 71
rect -1573 21 -1453 37
rect -1395 71 -1275 109
rect -1395 37 -1379 71
rect -1291 37 -1275 71
rect -1395 21 -1275 37
rect -1217 71 -1097 109
rect -1217 37 -1201 71
rect -1113 37 -1097 71
rect -1217 21 -1097 37
rect -1039 71 -919 109
rect -1039 37 -1023 71
rect -935 37 -919 71
rect -1039 21 -919 37
rect -861 71 -741 109
rect -861 37 -845 71
rect -757 37 -741 71
rect -861 21 -741 37
rect -683 71 -563 109
rect -683 37 -667 71
rect -579 37 -563 71
rect -683 21 -563 37
rect -505 71 -385 109
rect -505 37 -489 71
rect -401 37 -385 71
rect -505 21 -385 37
rect -327 71 -207 109
rect -327 37 -311 71
rect -223 37 -207 71
rect -327 21 -207 37
rect -149 71 -29 109
rect -149 37 -133 71
rect -45 37 -29 71
rect -149 21 -29 37
rect 29 71 149 109
rect 29 37 45 71
rect 133 37 149 71
rect 29 21 149 37
rect 207 71 327 109
rect 207 37 223 71
rect 311 37 327 71
rect 207 21 327 37
rect 385 71 505 109
rect 385 37 401 71
rect 489 37 505 71
rect 385 21 505 37
rect 563 71 683 109
rect 563 37 579 71
rect 667 37 683 71
rect 563 21 683 37
rect 741 71 861 109
rect 741 37 757 71
rect 845 37 861 71
rect 741 21 861 37
rect 919 71 1039 109
rect 919 37 935 71
rect 1023 37 1039 71
rect 919 21 1039 37
rect 1097 71 1217 109
rect 1097 37 1113 71
rect 1201 37 1217 71
rect 1097 21 1217 37
rect 1275 71 1395 109
rect 1275 37 1291 71
rect 1379 37 1395 71
rect 1275 21 1395 37
rect 1453 71 1573 109
rect 1453 37 1469 71
rect 1557 37 1573 71
rect 1453 21 1573 37
rect 1631 71 1751 109
rect 1631 37 1647 71
rect 1735 37 1751 71
rect 1631 21 1751 37
rect -1751 -37 -1631 -21
rect -1751 -71 -1735 -37
rect -1647 -71 -1631 -37
rect -1751 -109 -1631 -71
rect -1573 -37 -1453 -21
rect -1573 -71 -1557 -37
rect -1469 -71 -1453 -37
rect -1573 -109 -1453 -71
rect -1395 -37 -1275 -21
rect -1395 -71 -1379 -37
rect -1291 -71 -1275 -37
rect -1395 -109 -1275 -71
rect -1217 -37 -1097 -21
rect -1217 -71 -1201 -37
rect -1113 -71 -1097 -37
rect -1217 -109 -1097 -71
rect -1039 -37 -919 -21
rect -1039 -71 -1023 -37
rect -935 -71 -919 -37
rect -1039 -109 -919 -71
rect -861 -37 -741 -21
rect -861 -71 -845 -37
rect -757 -71 -741 -37
rect -861 -109 -741 -71
rect -683 -37 -563 -21
rect -683 -71 -667 -37
rect -579 -71 -563 -37
rect -683 -109 -563 -71
rect -505 -37 -385 -21
rect -505 -71 -489 -37
rect -401 -71 -385 -37
rect -505 -109 -385 -71
rect -327 -37 -207 -21
rect -327 -71 -311 -37
rect -223 -71 -207 -37
rect -327 -109 -207 -71
rect -149 -37 -29 -21
rect -149 -71 -133 -37
rect -45 -71 -29 -37
rect -149 -109 -29 -71
rect 29 -37 149 -21
rect 29 -71 45 -37
rect 133 -71 149 -37
rect 29 -109 149 -71
rect 207 -37 327 -21
rect 207 -71 223 -37
rect 311 -71 327 -37
rect 207 -109 327 -71
rect 385 -37 505 -21
rect 385 -71 401 -37
rect 489 -71 505 -37
rect 385 -109 505 -71
rect 563 -37 683 -21
rect 563 -71 579 -37
rect 667 -71 683 -37
rect 563 -109 683 -71
rect 741 -37 861 -21
rect 741 -71 757 -37
rect 845 -71 861 -37
rect 741 -109 861 -71
rect 919 -37 1039 -21
rect 919 -71 935 -37
rect 1023 -71 1039 -37
rect 919 -109 1039 -71
rect 1097 -37 1217 -21
rect 1097 -71 1113 -37
rect 1201 -71 1217 -37
rect 1097 -109 1217 -71
rect 1275 -37 1395 -21
rect 1275 -71 1291 -37
rect 1379 -71 1395 -37
rect 1275 -109 1395 -71
rect 1453 -37 1573 -21
rect 1453 -71 1469 -37
rect 1557 -71 1573 -37
rect 1453 -109 1573 -71
rect 1631 -37 1751 -21
rect 1631 -71 1647 -37
rect 1735 -71 1751 -37
rect 1631 -109 1751 -71
rect -1751 -1347 -1631 -1309
rect -1751 -1381 -1735 -1347
rect -1647 -1381 -1631 -1347
rect -1751 -1397 -1631 -1381
rect -1573 -1347 -1453 -1309
rect -1573 -1381 -1557 -1347
rect -1469 -1381 -1453 -1347
rect -1573 -1397 -1453 -1381
rect -1395 -1347 -1275 -1309
rect -1395 -1381 -1379 -1347
rect -1291 -1381 -1275 -1347
rect -1395 -1397 -1275 -1381
rect -1217 -1347 -1097 -1309
rect -1217 -1381 -1201 -1347
rect -1113 -1381 -1097 -1347
rect -1217 -1397 -1097 -1381
rect -1039 -1347 -919 -1309
rect -1039 -1381 -1023 -1347
rect -935 -1381 -919 -1347
rect -1039 -1397 -919 -1381
rect -861 -1347 -741 -1309
rect -861 -1381 -845 -1347
rect -757 -1381 -741 -1347
rect -861 -1397 -741 -1381
rect -683 -1347 -563 -1309
rect -683 -1381 -667 -1347
rect -579 -1381 -563 -1347
rect -683 -1397 -563 -1381
rect -505 -1347 -385 -1309
rect -505 -1381 -489 -1347
rect -401 -1381 -385 -1347
rect -505 -1397 -385 -1381
rect -327 -1347 -207 -1309
rect -327 -1381 -311 -1347
rect -223 -1381 -207 -1347
rect -327 -1397 -207 -1381
rect -149 -1347 -29 -1309
rect -149 -1381 -133 -1347
rect -45 -1381 -29 -1347
rect -149 -1397 -29 -1381
rect 29 -1347 149 -1309
rect 29 -1381 45 -1347
rect 133 -1381 149 -1347
rect 29 -1397 149 -1381
rect 207 -1347 327 -1309
rect 207 -1381 223 -1347
rect 311 -1381 327 -1347
rect 207 -1397 327 -1381
rect 385 -1347 505 -1309
rect 385 -1381 401 -1347
rect 489 -1381 505 -1347
rect 385 -1397 505 -1381
rect 563 -1347 683 -1309
rect 563 -1381 579 -1347
rect 667 -1381 683 -1347
rect 563 -1397 683 -1381
rect 741 -1347 861 -1309
rect 741 -1381 757 -1347
rect 845 -1381 861 -1347
rect 741 -1397 861 -1381
rect 919 -1347 1039 -1309
rect 919 -1381 935 -1347
rect 1023 -1381 1039 -1347
rect 919 -1397 1039 -1381
rect 1097 -1347 1217 -1309
rect 1097 -1381 1113 -1347
rect 1201 -1381 1217 -1347
rect 1097 -1397 1217 -1381
rect 1275 -1347 1395 -1309
rect 1275 -1381 1291 -1347
rect 1379 -1381 1395 -1347
rect 1275 -1397 1395 -1381
rect 1453 -1347 1573 -1309
rect 1453 -1381 1469 -1347
rect 1557 -1381 1573 -1347
rect 1453 -1397 1573 -1381
rect 1631 -1347 1751 -1309
rect 1631 -1381 1647 -1347
rect 1735 -1381 1751 -1347
rect 1631 -1397 1751 -1381
<< polycont >>
rect -1735 1347 -1647 1381
rect -1557 1347 -1469 1381
rect -1379 1347 -1291 1381
rect -1201 1347 -1113 1381
rect -1023 1347 -935 1381
rect -845 1347 -757 1381
rect -667 1347 -579 1381
rect -489 1347 -401 1381
rect -311 1347 -223 1381
rect -133 1347 -45 1381
rect 45 1347 133 1381
rect 223 1347 311 1381
rect 401 1347 489 1381
rect 579 1347 667 1381
rect 757 1347 845 1381
rect 935 1347 1023 1381
rect 1113 1347 1201 1381
rect 1291 1347 1379 1381
rect 1469 1347 1557 1381
rect 1647 1347 1735 1381
rect -1735 37 -1647 71
rect -1557 37 -1469 71
rect -1379 37 -1291 71
rect -1201 37 -1113 71
rect -1023 37 -935 71
rect -845 37 -757 71
rect -667 37 -579 71
rect -489 37 -401 71
rect -311 37 -223 71
rect -133 37 -45 71
rect 45 37 133 71
rect 223 37 311 71
rect 401 37 489 71
rect 579 37 667 71
rect 757 37 845 71
rect 935 37 1023 71
rect 1113 37 1201 71
rect 1291 37 1379 71
rect 1469 37 1557 71
rect 1647 37 1735 71
rect -1735 -71 -1647 -37
rect -1557 -71 -1469 -37
rect -1379 -71 -1291 -37
rect -1201 -71 -1113 -37
rect -1023 -71 -935 -37
rect -845 -71 -757 -37
rect -667 -71 -579 -37
rect -489 -71 -401 -37
rect -311 -71 -223 -37
rect -133 -71 -45 -37
rect 45 -71 133 -37
rect 223 -71 311 -37
rect 401 -71 489 -37
rect 579 -71 667 -37
rect 757 -71 845 -37
rect 935 -71 1023 -37
rect 1113 -71 1201 -37
rect 1291 -71 1379 -37
rect 1469 -71 1557 -37
rect 1647 -71 1735 -37
rect -1735 -1381 -1647 -1347
rect -1557 -1381 -1469 -1347
rect -1379 -1381 -1291 -1347
rect -1201 -1381 -1113 -1347
rect -1023 -1381 -935 -1347
rect -845 -1381 -757 -1347
rect -667 -1381 -579 -1347
rect -489 -1381 -401 -1347
rect -311 -1381 -223 -1347
rect -133 -1381 -45 -1347
rect 45 -1381 133 -1347
rect 223 -1381 311 -1347
rect 401 -1381 489 -1347
rect 579 -1381 667 -1347
rect 757 -1381 845 -1347
rect 935 -1381 1023 -1347
rect 1113 -1381 1201 -1347
rect 1291 -1381 1379 -1347
rect 1469 -1381 1557 -1347
rect 1647 -1381 1735 -1347
<< locali >>
rect -1911 1449 -1815 1483
rect 1815 1449 1911 1483
rect -1911 1387 -1877 1449
rect 1877 1387 1911 1449
rect -1751 1347 -1735 1381
rect -1647 1347 -1631 1381
rect -1573 1347 -1557 1381
rect -1469 1347 -1453 1381
rect -1395 1347 -1379 1381
rect -1291 1347 -1275 1381
rect -1217 1347 -1201 1381
rect -1113 1347 -1097 1381
rect -1039 1347 -1023 1381
rect -935 1347 -919 1381
rect -861 1347 -845 1381
rect -757 1347 -741 1381
rect -683 1347 -667 1381
rect -579 1347 -563 1381
rect -505 1347 -489 1381
rect -401 1347 -385 1381
rect -327 1347 -311 1381
rect -223 1347 -207 1381
rect -149 1347 -133 1381
rect -45 1347 -29 1381
rect 29 1347 45 1381
rect 133 1347 149 1381
rect 207 1347 223 1381
rect 311 1347 327 1381
rect 385 1347 401 1381
rect 489 1347 505 1381
rect 563 1347 579 1381
rect 667 1347 683 1381
rect 741 1347 757 1381
rect 845 1347 861 1381
rect 919 1347 935 1381
rect 1023 1347 1039 1381
rect 1097 1347 1113 1381
rect 1201 1347 1217 1381
rect 1275 1347 1291 1381
rect 1379 1347 1395 1381
rect 1453 1347 1469 1381
rect 1557 1347 1573 1381
rect 1631 1347 1647 1381
rect 1735 1347 1751 1381
rect -1797 1297 -1763 1313
rect -1797 105 -1763 121
rect -1619 1297 -1585 1313
rect -1619 105 -1585 121
rect -1441 1297 -1407 1313
rect -1441 105 -1407 121
rect -1263 1297 -1229 1313
rect -1263 105 -1229 121
rect -1085 1297 -1051 1313
rect -1085 105 -1051 121
rect -907 1297 -873 1313
rect -907 105 -873 121
rect -729 1297 -695 1313
rect -729 105 -695 121
rect -551 1297 -517 1313
rect -551 105 -517 121
rect -373 1297 -339 1313
rect -373 105 -339 121
rect -195 1297 -161 1313
rect -195 105 -161 121
rect -17 1297 17 1313
rect -17 105 17 121
rect 161 1297 195 1313
rect 161 105 195 121
rect 339 1297 373 1313
rect 339 105 373 121
rect 517 1297 551 1313
rect 517 105 551 121
rect 695 1297 729 1313
rect 695 105 729 121
rect 873 1297 907 1313
rect 873 105 907 121
rect 1051 1297 1085 1313
rect 1051 105 1085 121
rect 1229 1297 1263 1313
rect 1229 105 1263 121
rect 1407 1297 1441 1313
rect 1407 105 1441 121
rect 1585 1297 1619 1313
rect 1585 105 1619 121
rect 1763 1297 1797 1313
rect 1763 105 1797 121
rect -1751 37 -1735 71
rect -1647 37 -1631 71
rect -1573 37 -1557 71
rect -1469 37 -1453 71
rect -1395 37 -1379 71
rect -1291 37 -1275 71
rect -1217 37 -1201 71
rect -1113 37 -1097 71
rect -1039 37 -1023 71
rect -935 37 -919 71
rect -861 37 -845 71
rect -757 37 -741 71
rect -683 37 -667 71
rect -579 37 -563 71
rect -505 37 -489 71
rect -401 37 -385 71
rect -327 37 -311 71
rect -223 37 -207 71
rect -149 37 -133 71
rect -45 37 -29 71
rect 29 37 45 71
rect 133 37 149 71
rect 207 37 223 71
rect 311 37 327 71
rect 385 37 401 71
rect 489 37 505 71
rect 563 37 579 71
rect 667 37 683 71
rect 741 37 757 71
rect 845 37 861 71
rect 919 37 935 71
rect 1023 37 1039 71
rect 1097 37 1113 71
rect 1201 37 1217 71
rect 1275 37 1291 71
rect 1379 37 1395 71
rect 1453 37 1469 71
rect 1557 37 1573 71
rect 1631 37 1647 71
rect 1735 37 1751 71
rect -1751 -71 -1735 -37
rect -1647 -71 -1631 -37
rect -1573 -71 -1557 -37
rect -1469 -71 -1453 -37
rect -1395 -71 -1379 -37
rect -1291 -71 -1275 -37
rect -1217 -71 -1201 -37
rect -1113 -71 -1097 -37
rect -1039 -71 -1023 -37
rect -935 -71 -919 -37
rect -861 -71 -845 -37
rect -757 -71 -741 -37
rect -683 -71 -667 -37
rect -579 -71 -563 -37
rect -505 -71 -489 -37
rect -401 -71 -385 -37
rect -327 -71 -311 -37
rect -223 -71 -207 -37
rect -149 -71 -133 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 133 -71 149 -37
rect 207 -71 223 -37
rect 311 -71 327 -37
rect 385 -71 401 -37
rect 489 -71 505 -37
rect 563 -71 579 -37
rect 667 -71 683 -37
rect 741 -71 757 -37
rect 845 -71 861 -37
rect 919 -71 935 -37
rect 1023 -71 1039 -37
rect 1097 -71 1113 -37
rect 1201 -71 1217 -37
rect 1275 -71 1291 -37
rect 1379 -71 1395 -37
rect 1453 -71 1469 -37
rect 1557 -71 1573 -37
rect 1631 -71 1647 -37
rect 1735 -71 1751 -37
rect -1797 -121 -1763 -105
rect -1797 -1313 -1763 -1297
rect -1619 -121 -1585 -105
rect -1619 -1313 -1585 -1297
rect -1441 -121 -1407 -105
rect -1441 -1313 -1407 -1297
rect -1263 -121 -1229 -105
rect -1263 -1313 -1229 -1297
rect -1085 -121 -1051 -105
rect -1085 -1313 -1051 -1297
rect -907 -121 -873 -105
rect -907 -1313 -873 -1297
rect -729 -121 -695 -105
rect -729 -1313 -695 -1297
rect -551 -121 -517 -105
rect -551 -1313 -517 -1297
rect -373 -121 -339 -105
rect -373 -1313 -339 -1297
rect -195 -121 -161 -105
rect -195 -1313 -161 -1297
rect -17 -121 17 -105
rect -17 -1313 17 -1297
rect 161 -121 195 -105
rect 161 -1313 195 -1297
rect 339 -121 373 -105
rect 339 -1313 373 -1297
rect 517 -121 551 -105
rect 517 -1313 551 -1297
rect 695 -121 729 -105
rect 695 -1313 729 -1297
rect 873 -121 907 -105
rect 873 -1313 907 -1297
rect 1051 -121 1085 -105
rect 1051 -1313 1085 -1297
rect 1229 -121 1263 -105
rect 1229 -1313 1263 -1297
rect 1407 -121 1441 -105
rect 1407 -1313 1441 -1297
rect 1585 -121 1619 -105
rect 1585 -1313 1619 -1297
rect 1763 -121 1797 -105
rect 1763 -1313 1797 -1297
rect -1751 -1381 -1735 -1347
rect -1647 -1381 -1631 -1347
rect -1573 -1381 -1557 -1347
rect -1469 -1381 -1453 -1347
rect -1395 -1381 -1379 -1347
rect -1291 -1381 -1275 -1347
rect -1217 -1381 -1201 -1347
rect -1113 -1381 -1097 -1347
rect -1039 -1381 -1023 -1347
rect -935 -1381 -919 -1347
rect -861 -1381 -845 -1347
rect -757 -1381 -741 -1347
rect -683 -1381 -667 -1347
rect -579 -1381 -563 -1347
rect -505 -1381 -489 -1347
rect -401 -1381 -385 -1347
rect -327 -1381 -311 -1347
rect -223 -1381 -207 -1347
rect -149 -1381 -133 -1347
rect -45 -1381 -29 -1347
rect 29 -1381 45 -1347
rect 133 -1381 149 -1347
rect 207 -1381 223 -1347
rect 311 -1381 327 -1347
rect 385 -1381 401 -1347
rect 489 -1381 505 -1347
rect 563 -1381 579 -1347
rect 667 -1381 683 -1347
rect 741 -1381 757 -1347
rect 845 -1381 861 -1347
rect 919 -1381 935 -1347
rect 1023 -1381 1039 -1347
rect 1097 -1381 1113 -1347
rect 1201 -1381 1217 -1347
rect 1275 -1381 1291 -1347
rect 1379 -1381 1395 -1347
rect 1453 -1381 1469 -1347
rect 1557 -1381 1573 -1347
rect 1631 -1381 1647 -1347
rect 1735 -1381 1751 -1347
rect -1911 -1449 -1877 -1387
rect 1877 -1449 1911 -1387
rect -1911 -1483 -1815 -1449
rect 1815 -1483 1911 -1449
<< viali >>
rect -1735 1347 -1647 1381
rect -1557 1347 -1469 1381
rect -1379 1347 -1291 1381
rect -1201 1347 -1113 1381
rect -1023 1347 -935 1381
rect -845 1347 -757 1381
rect -667 1347 -579 1381
rect -489 1347 -401 1381
rect -311 1347 -223 1381
rect -133 1347 -45 1381
rect 45 1347 133 1381
rect 223 1347 311 1381
rect 401 1347 489 1381
rect 579 1347 667 1381
rect 757 1347 845 1381
rect 935 1347 1023 1381
rect 1113 1347 1201 1381
rect 1291 1347 1379 1381
rect 1469 1347 1557 1381
rect 1647 1347 1735 1381
rect -1797 121 -1763 1297
rect -1619 121 -1585 1297
rect -1441 121 -1407 1297
rect -1263 121 -1229 1297
rect -1085 121 -1051 1297
rect -907 121 -873 1297
rect -729 121 -695 1297
rect -551 121 -517 1297
rect -373 121 -339 1297
rect -195 121 -161 1297
rect -17 121 17 1297
rect 161 121 195 1297
rect 339 121 373 1297
rect 517 121 551 1297
rect 695 121 729 1297
rect 873 121 907 1297
rect 1051 121 1085 1297
rect 1229 121 1263 1297
rect 1407 121 1441 1297
rect 1585 121 1619 1297
rect 1763 121 1797 1297
rect -1735 37 -1647 71
rect -1557 37 -1469 71
rect -1379 37 -1291 71
rect -1201 37 -1113 71
rect -1023 37 -935 71
rect -845 37 -757 71
rect -667 37 -579 71
rect -489 37 -401 71
rect -311 37 -223 71
rect -133 37 -45 71
rect 45 37 133 71
rect 223 37 311 71
rect 401 37 489 71
rect 579 37 667 71
rect 757 37 845 71
rect 935 37 1023 71
rect 1113 37 1201 71
rect 1291 37 1379 71
rect 1469 37 1557 71
rect 1647 37 1735 71
rect -1735 -71 -1647 -37
rect -1557 -71 -1469 -37
rect -1379 -71 -1291 -37
rect -1201 -71 -1113 -37
rect -1023 -71 -935 -37
rect -845 -71 -757 -37
rect -667 -71 -579 -37
rect -489 -71 -401 -37
rect -311 -71 -223 -37
rect -133 -71 -45 -37
rect 45 -71 133 -37
rect 223 -71 311 -37
rect 401 -71 489 -37
rect 579 -71 667 -37
rect 757 -71 845 -37
rect 935 -71 1023 -37
rect 1113 -71 1201 -37
rect 1291 -71 1379 -37
rect 1469 -71 1557 -37
rect 1647 -71 1735 -37
rect -1797 -1297 -1763 -121
rect -1619 -1297 -1585 -121
rect -1441 -1297 -1407 -121
rect -1263 -1297 -1229 -121
rect -1085 -1297 -1051 -121
rect -907 -1297 -873 -121
rect -729 -1297 -695 -121
rect -551 -1297 -517 -121
rect -373 -1297 -339 -121
rect -195 -1297 -161 -121
rect -17 -1297 17 -121
rect 161 -1297 195 -121
rect 339 -1297 373 -121
rect 517 -1297 551 -121
rect 695 -1297 729 -121
rect 873 -1297 907 -121
rect 1051 -1297 1085 -121
rect 1229 -1297 1263 -121
rect 1407 -1297 1441 -121
rect 1585 -1297 1619 -121
rect 1763 -1297 1797 -121
rect -1735 -1381 -1647 -1347
rect -1557 -1381 -1469 -1347
rect -1379 -1381 -1291 -1347
rect -1201 -1381 -1113 -1347
rect -1023 -1381 -935 -1347
rect -845 -1381 -757 -1347
rect -667 -1381 -579 -1347
rect -489 -1381 -401 -1347
rect -311 -1381 -223 -1347
rect -133 -1381 -45 -1347
rect 45 -1381 133 -1347
rect 223 -1381 311 -1347
rect 401 -1381 489 -1347
rect 579 -1381 667 -1347
rect 757 -1381 845 -1347
rect 935 -1381 1023 -1347
rect 1113 -1381 1201 -1347
rect 1291 -1381 1379 -1347
rect 1469 -1381 1557 -1347
rect 1647 -1381 1735 -1347
<< metal1 >>
rect -1747 1381 -1635 1387
rect -1747 1347 -1735 1381
rect -1647 1347 -1635 1381
rect -1747 1341 -1635 1347
rect -1569 1381 -1457 1387
rect -1569 1347 -1557 1381
rect -1469 1347 -1457 1381
rect -1569 1341 -1457 1347
rect -1391 1381 -1279 1387
rect -1391 1347 -1379 1381
rect -1291 1347 -1279 1381
rect -1391 1341 -1279 1347
rect -1213 1381 -1101 1387
rect -1213 1347 -1201 1381
rect -1113 1347 -1101 1381
rect -1213 1341 -1101 1347
rect -1035 1381 -923 1387
rect -1035 1347 -1023 1381
rect -935 1347 -923 1381
rect -1035 1341 -923 1347
rect -857 1381 -745 1387
rect -857 1347 -845 1381
rect -757 1347 -745 1381
rect -857 1341 -745 1347
rect -679 1381 -567 1387
rect -679 1347 -667 1381
rect -579 1347 -567 1381
rect -679 1341 -567 1347
rect -501 1381 -389 1387
rect -501 1347 -489 1381
rect -401 1347 -389 1381
rect -501 1341 -389 1347
rect -323 1381 -211 1387
rect -323 1347 -311 1381
rect -223 1347 -211 1381
rect -323 1341 -211 1347
rect -145 1381 -33 1387
rect -145 1347 -133 1381
rect -45 1347 -33 1381
rect -145 1341 -33 1347
rect 33 1381 145 1387
rect 33 1347 45 1381
rect 133 1347 145 1381
rect 33 1341 145 1347
rect 211 1381 323 1387
rect 211 1347 223 1381
rect 311 1347 323 1381
rect 211 1341 323 1347
rect 389 1381 501 1387
rect 389 1347 401 1381
rect 489 1347 501 1381
rect 389 1341 501 1347
rect 567 1381 679 1387
rect 567 1347 579 1381
rect 667 1347 679 1381
rect 567 1341 679 1347
rect 745 1381 857 1387
rect 745 1347 757 1381
rect 845 1347 857 1381
rect 745 1341 857 1347
rect 923 1381 1035 1387
rect 923 1347 935 1381
rect 1023 1347 1035 1381
rect 923 1341 1035 1347
rect 1101 1381 1213 1387
rect 1101 1347 1113 1381
rect 1201 1347 1213 1381
rect 1101 1341 1213 1347
rect 1279 1381 1391 1387
rect 1279 1347 1291 1381
rect 1379 1347 1391 1381
rect 1279 1341 1391 1347
rect 1457 1381 1569 1387
rect 1457 1347 1469 1381
rect 1557 1347 1569 1381
rect 1457 1341 1569 1347
rect 1635 1381 1747 1387
rect 1635 1347 1647 1381
rect 1735 1347 1747 1381
rect 1635 1341 1747 1347
rect -1803 1297 -1757 1309
rect -1803 121 -1797 1297
rect -1763 121 -1757 1297
rect -1803 109 -1757 121
rect -1625 1297 -1579 1309
rect -1625 121 -1619 1297
rect -1585 121 -1579 1297
rect -1625 109 -1579 121
rect -1447 1297 -1401 1309
rect -1447 121 -1441 1297
rect -1407 121 -1401 1297
rect -1447 109 -1401 121
rect -1269 1297 -1223 1309
rect -1269 121 -1263 1297
rect -1229 121 -1223 1297
rect -1269 109 -1223 121
rect -1091 1297 -1045 1309
rect -1091 121 -1085 1297
rect -1051 121 -1045 1297
rect -1091 109 -1045 121
rect -913 1297 -867 1309
rect -913 121 -907 1297
rect -873 121 -867 1297
rect -913 109 -867 121
rect -735 1297 -689 1309
rect -735 121 -729 1297
rect -695 121 -689 1297
rect -735 109 -689 121
rect -557 1297 -511 1309
rect -557 121 -551 1297
rect -517 121 -511 1297
rect -557 109 -511 121
rect -379 1297 -333 1309
rect -379 121 -373 1297
rect -339 121 -333 1297
rect -379 109 -333 121
rect -201 1297 -155 1309
rect -201 121 -195 1297
rect -161 121 -155 1297
rect -201 109 -155 121
rect -23 1297 23 1309
rect -23 121 -17 1297
rect 17 121 23 1297
rect -23 109 23 121
rect 155 1297 201 1309
rect 155 121 161 1297
rect 195 121 201 1297
rect 155 109 201 121
rect 333 1297 379 1309
rect 333 121 339 1297
rect 373 121 379 1297
rect 333 109 379 121
rect 511 1297 557 1309
rect 511 121 517 1297
rect 551 121 557 1297
rect 511 109 557 121
rect 689 1297 735 1309
rect 689 121 695 1297
rect 729 121 735 1297
rect 689 109 735 121
rect 867 1297 913 1309
rect 867 121 873 1297
rect 907 121 913 1297
rect 867 109 913 121
rect 1045 1297 1091 1309
rect 1045 121 1051 1297
rect 1085 121 1091 1297
rect 1045 109 1091 121
rect 1223 1297 1269 1309
rect 1223 121 1229 1297
rect 1263 121 1269 1297
rect 1223 109 1269 121
rect 1401 1297 1447 1309
rect 1401 121 1407 1297
rect 1441 121 1447 1297
rect 1401 109 1447 121
rect 1579 1297 1625 1309
rect 1579 121 1585 1297
rect 1619 121 1625 1297
rect 1579 109 1625 121
rect 1757 1297 1803 1309
rect 1757 121 1763 1297
rect 1797 121 1803 1297
rect 1757 109 1803 121
rect -1747 71 -1635 77
rect -1747 37 -1735 71
rect -1647 37 -1635 71
rect -1747 31 -1635 37
rect -1569 71 -1457 77
rect -1569 37 -1557 71
rect -1469 37 -1457 71
rect -1569 31 -1457 37
rect -1391 71 -1279 77
rect -1391 37 -1379 71
rect -1291 37 -1279 71
rect -1391 31 -1279 37
rect -1213 71 -1101 77
rect -1213 37 -1201 71
rect -1113 37 -1101 71
rect -1213 31 -1101 37
rect -1035 71 -923 77
rect -1035 37 -1023 71
rect -935 37 -923 71
rect -1035 31 -923 37
rect -857 71 -745 77
rect -857 37 -845 71
rect -757 37 -745 71
rect -857 31 -745 37
rect -679 71 -567 77
rect -679 37 -667 71
rect -579 37 -567 71
rect -679 31 -567 37
rect -501 71 -389 77
rect -501 37 -489 71
rect -401 37 -389 71
rect -501 31 -389 37
rect -323 71 -211 77
rect -323 37 -311 71
rect -223 37 -211 71
rect -323 31 -211 37
rect -145 71 -33 77
rect -145 37 -133 71
rect -45 37 -33 71
rect -145 31 -33 37
rect 33 71 145 77
rect 33 37 45 71
rect 133 37 145 71
rect 33 31 145 37
rect 211 71 323 77
rect 211 37 223 71
rect 311 37 323 71
rect 211 31 323 37
rect 389 71 501 77
rect 389 37 401 71
rect 489 37 501 71
rect 389 31 501 37
rect 567 71 679 77
rect 567 37 579 71
rect 667 37 679 71
rect 567 31 679 37
rect 745 71 857 77
rect 745 37 757 71
rect 845 37 857 71
rect 745 31 857 37
rect 923 71 1035 77
rect 923 37 935 71
rect 1023 37 1035 71
rect 923 31 1035 37
rect 1101 71 1213 77
rect 1101 37 1113 71
rect 1201 37 1213 71
rect 1101 31 1213 37
rect 1279 71 1391 77
rect 1279 37 1291 71
rect 1379 37 1391 71
rect 1279 31 1391 37
rect 1457 71 1569 77
rect 1457 37 1469 71
rect 1557 37 1569 71
rect 1457 31 1569 37
rect 1635 71 1747 77
rect 1635 37 1647 71
rect 1735 37 1747 71
rect 1635 31 1747 37
rect -1747 -37 -1635 -31
rect -1747 -71 -1735 -37
rect -1647 -71 -1635 -37
rect -1747 -77 -1635 -71
rect -1569 -37 -1457 -31
rect -1569 -71 -1557 -37
rect -1469 -71 -1457 -37
rect -1569 -77 -1457 -71
rect -1391 -37 -1279 -31
rect -1391 -71 -1379 -37
rect -1291 -71 -1279 -37
rect -1391 -77 -1279 -71
rect -1213 -37 -1101 -31
rect -1213 -71 -1201 -37
rect -1113 -71 -1101 -37
rect -1213 -77 -1101 -71
rect -1035 -37 -923 -31
rect -1035 -71 -1023 -37
rect -935 -71 -923 -37
rect -1035 -77 -923 -71
rect -857 -37 -745 -31
rect -857 -71 -845 -37
rect -757 -71 -745 -37
rect -857 -77 -745 -71
rect -679 -37 -567 -31
rect -679 -71 -667 -37
rect -579 -71 -567 -37
rect -679 -77 -567 -71
rect -501 -37 -389 -31
rect -501 -71 -489 -37
rect -401 -71 -389 -37
rect -501 -77 -389 -71
rect -323 -37 -211 -31
rect -323 -71 -311 -37
rect -223 -71 -211 -37
rect -323 -77 -211 -71
rect -145 -37 -33 -31
rect -145 -71 -133 -37
rect -45 -71 -33 -37
rect -145 -77 -33 -71
rect 33 -37 145 -31
rect 33 -71 45 -37
rect 133 -71 145 -37
rect 33 -77 145 -71
rect 211 -37 323 -31
rect 211 -71 223 -37
rect 311 -71 323 -37
rect 211 -77 323 -71
rect 389 -37 501 -31
rect 389 -71 401 -37
rect 489 -71 501 -37
rect 389 -77 501 -71
rect 567 -37 679 -31
rect 567 -71 579 -37
rect 667 -71 679 -37
rect 567 -77 679 -71
rect 745 -37 857 -31
rect 745 -71 757 -37
rect 845 -71 857 -37
rect 745 -77 857 -71
rect 923 -37 1035 -31
rect 923 -71 935 -37
rect 1023 -71 1035 -37
rect 923 -77 1035 -71
rect 1101 -37 1213 -31
rect 1101 -71 1113 -37
rect 1201 -71 1213 -37
rect 1101 -77 1213 -71
rect 1279 -37 1391 -31
rect 1279 -71 1291 -37
rect 1379 -71 1391 -37
rect 1279 -77 1391 -71
rect 1457 -37 1569 -31
rect 1457 -71 1469 -37
rect 1557 -71 1569 -37
rect 1457 -77 1569 -71
rect 1635 -37 1747 -31
rect 1635 -71 1647 -37
rect 1735 -71 1747 -37
rect 1635 -77 1747 -71
rect -1803 -121 -1757 -109
rect -1803 -1297 -1797 -121
rect -1763 -1297 -1757 -121
rect -1803 -1309 -1757 -1297
rect -1625 -121 -1579 -109
rect -1625 -1297 -1619 -121
rect -1585 -1297 -1579 -121
rect -1625 -1309 -1579 -1297
rect -1447 -121 -1401 -109
rect -1447 -1297 -1441 -121
rect -1407 -1297 -1401 -121
rect -1447 -1309 -1401 -1297
rect -1269 -121 -1223 -109
rect -1269 -1297 -1263 -121
rect -1229 -1297 -1223 -121
rect -1269 -1309 -1223 -1297
rect -1091 -121 -1045 -109
rect -1091 -1297 -1085 -121
rect -1051 -1297 -1045 -121
rect -1091 -1309 -1045 -1297
rect -913 -121 -867 -109
rect -913 -1297 -907 -121
rect -873 -1297 -867 -121
rect -913 -1309 -867 -1297
rect -735 -121 -689 -109
rect -735 -1297 -729 -121
rect -695 -1297 -689 -121
rect -735 -1309 -689 -1297
rect -557 -121 -511 -109
rect -557 -1297 -551 -121
rect -517 -1297 -511 -121
rect -557 -1309 -511 -1297
rect -379 -121 -333 -109
rect -379 -1297 -373 -121
rect -339 -1297 -333 -121
rect -379 -1309 -333 -1297
rect -201 -121 -155 -109
rect -201 -1297 -195 -121
rect -161 -1297 -155 -121
rect -201 -1309 -155 -1297
rect -23 -121 23 -109
rect -23 -1297 -17 -121
rect 17 -1297 23 -121
rect -23 -1309 23 -1297
rect 155 -121 201 -109
rect 155 -1297 161 -121
rect 195 -1297 201 -121
rect 155 -1309 201 -1297
rect 333 -121 379 -109
rect 333 -1297 339 -121
rect 373 -1297 379 -121
rect 333 -1309 379 -1297
rect 511 -121 557 -109
rect 511 -1297 517 -121
rect 551 -1297 557 -121
rect 511 -1309 557 -1297
rect 689 -121 735 -109
rect 689 -1297 695 -121
rect 729 -1297 735 -121
rect 689 -1309 735 -1297
rect 867 -121 913 -109
rect 867 -1297 873 -121
rect 907 -1297 913 -121
rect 867 -1309 913 -1297
rect 1045 -121 1091 -109
rect 1045 -1297 1051 -121
rect 1085 -1297 1091 -121
rect 1045 -1309 1091 -1297
rect 1223 -121 1269 -109
rect 1223 -1297 1229 -121
rect 1263 -1297 1269 -121
rect 1223 -1309 1269 -1297
rect 1401 -121 1447 -109
rect 1401 -1297 1407 -121
rect 1441 -1297 1447 -121
rect 1401 -1309 1447 -1297
rect 1579 -121 1625 -109
rect 1579 -1297 1585 -121
rect 1619 -1297 1625 -121
rect 1579 -1309 1625 -1297
rect 1757 -121 1803 -109
rect 1757 -1297 1763 -121
rect 1797 -1297 1803 -121
rect 1757 -1309 1803 -1297
rect -1747 -1347 -1635 -1341
rect -1747 -1381 -1735 -1347
rect -1647 -1381 -1635 -1347
rect -1747 -1387 -1635 -1381
rect -1569 -1347 -1457 -1341
rect -1569 -1381 -1557 -1347
rect -1469 -1381 -1457 -1347
rect -1569 -1387 -1457 -1381
rect -1391 -1347 -1279 -1341
rect -1391 -1381 -1379 -1347
rect -1291 -1381 -1279 -1347
rect -1391 -1387 -1279 -1381
rect -1213 -1347 -1101 -1341
rect -1213 -1381 -1201 -1347
rect -1113 -1381 -1101 -1347
rect -1213 -1387 -1101 -1381
rect -1035 -1347 -923 -1341
rect -1035 -1381 -1023 -1347
rect -935 -1381 -923 -1347
rect -1035 -1387 -923 -1381
rect -857 -1347 -745 -1341
rect -857 -1381 -845 -1347
rect -757 -1381 -745 -1347
rect -857 -1387 -745 -1381
rect -679 -1347 -567 -1341
rect -679 -1381 -667 -1347
rect -579 -1381 -567 -1347
rect -679 -1387 -567 -1381
rect -501 -1347 -389 -1341
rect -501 -1381 -489 -1347
rect -401 -1381 -389 -1347
rect -501 -1387 -389 -1381
rect -323 -1347 -211 -1341
rect -323 -1381 -311 -1347
rect -223 -1381 -211 -1347
rect -323 -1387 -211 -1381
rect -145 -1347 -33 -1341
rect -145 -1381 -133 -1347
rect -45 -1381 -33 -1347
rect -145 -1387 -33 -1381
rect 33 -1347 145 -1341
rect 33 -1381 45 -1347
rect 133 -1381 145 -1347
rect 33 -1387 145 -1381
rect 211 -1347 323 -1341
rect 211 -1381 223 -1347
rect 311 -1381 323 -1347
rect 211 -1387 323 -1381
rect 389 -1347 501 -1341
rect 389 -1381 401 -1347
rect 489 -1381 501 -1347
rect 389 -1387 501 -1381
rect 567 -1347 679 -1341
rect 567 -1381 579 -1347
rect 667 -1381 679 -1347
rect 567 -1387 679 -1381
rect 745 -1347 857 -1341
rect 745 -1381 757 -1347
rect 845 -1381 857 -1347
rect 745 -1387 857 -1381
rect 923 -1347 1035 -1341
rect 923 -1381 935 -1347
rect 1023 -1381 1035 -1347
rect 923 -1387 1035 -1381
rect 1101 -1347 1213 -1341
rect 1101 -1381 1113 -1347
rect 1201 -1381 1213 -1347
rect 1101 -1387 1213 -1381
rect 1279 -1347 1391 -1341
rect 1279 -1381 1291 -1347
rect 1379 -1381 1391 -1347
rect 1279 -1387 1391 -1381
rect 1457 -1347 1569 -1341
rect 1457 -1381 1469 -1347
rect 1557 -1381 1569 -1347
rect 1457 -1387 1569 -1381
rect 1635 -1347 1747 -1341
rect 1635 -1381 1647 -1347
rect 1735 -1381 1747 -1347
rect 1635 -1387 1747 -1381
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1894 -1466 1894 1466
string parameters w 6 l 0.6 m 2 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
