magic
tech sky130B
magscale 1 2
timestamp 1606424343
<< metal3 >>
rect -6924 1572 -3552 1600
rect -6924 -1572 -3636 1572
rect -3572 -1572 -3552 1572
rect -6924 -1600 -3552 -1572
rect -3432 1572 -60 1600
rect -3432 -1572 -144 1572
rect -80 -1572 -60 1572
rect -3432 -1600 -60 -1572
rect 60 1572 3432 1600
rect 60 -1572 3348 1572
rect 3412 -1572 3432 1572
rect 60 -1600 3432 -1572
rect 3552 1572 6924 1600
rect 3552 -1572 6840 1572
rect 6904 -1572 6924 1572
rect 3552 -1600 6924 -1572
<< via3 >>
rect -3636 -1572 -3572 1572
rect -144 -1572 -80 1572
rect 3348 -1572 3412 1572
rect 6840 -1572 6904 1572
<< mimcap >>
rect -6824 1460 -3824 1500
rect -6824 -1460 -6784 1460
rect -3864 -1460 -3824 1460
rect -6824 -1500 -3824 -1460
rect -3332 1460 -332 1500
rect -3332 -1460 -3292 1460
rect -372 -1460 -332 1460
rect -3332 -1500 -332 -1460
rect 160 1460 3160 1500
rect 160 -1460 200 1460
rect 3120 -1460 3160 1460
rect 160 -1500 3160 -1460
rect 3652 1460 6652 1500
rect 3652 -1460 3692 1460
rect 6612 -1460 6652 1460
rect 3652 -1500 6652 -1460
<< mimcapcontact >>
rect -6784 -1460 -3864 1460
rect -3292 -1460 -372 1460
rect 200 -1460 3120 1460
rect 3692 -1460 6612 1460
<< metal4 >>
rect -3652 1572 -3556 1588
rect -6785 1460 -3863 1461
rect -6785 -1460 -6784 1460
rect -3864 -1460 -3863 1460
rect -6785 -1461 -3863 -1460
rect -3652 -1572 -3636 1572
rect -3572 -1572 -3556 1572
rect -160 1572 -64 1588
rect -3293 1460 -371 1461
rect -3293 -1460 -3292 1460
rect -372 -1460 -371 1460
rect -3293 -1461 -371 -1460
rect -3652 -1588 -3556 -1572
rect -160 -1572 -144 1572
rect -80 -1572 -64 1572
rect 3332 1572 3428 1588
rect 199 1460 3121 1461
rect 199 -1460 200 1460
rect 3120 -1460 3121 1460
rect 199 -1461 3121 -1460
rect -160 -1588 -64 -1572
rect 3332 -1572 3348 1572
rect 3412 -1572 3428 1572
rect 6824 1572 6920 1588
rect 3691 1460 6613 1461
rect 3691 -1460 3692 1460
rect 6612 -1460 6613 1460
rect 3691 -1461 6613 -1460
rect 3332 -1588 3428 -1572
rect 6824 -1572 6840 1572
rect 6904 -1572 6920 1572
rect 6824 -1588 6920 -1572
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 3552 -1600 6752 1600
string parameters w 15.0 l 15.0 val 235.2 carea 1.00 cperi 0.17 nx 4 ny 1 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1
string library sky130
<< end >>
