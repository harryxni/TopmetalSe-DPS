magic
tech sky130B
magscale 1 2
timestamp 1662227450
<< nwell >>
rect -770 -3590 -1 -3240
rect 2520 -3590 3470 -3240
<< nmoslvt >>
rect 2590 -6880 2630 -5280
<< ndiff >>
rect 2520 -5310 2590 -5280
rect 2520 -6860 2530 -5310
rect 2570 -6860 2590 -5310
rect 2520 -6880 2590 -6860
rect 2630 -5310 2700 -5280
rect 2630 -6860 2650 -5310
rect 2690 -6860 2700 -5310
rect 2630 -6880 2700 -6860
<< ndiffc >>
rect 2530 -6860 2570 -5310
rect 2650 -6860 2690 -5310
<< poly >>
rect 2590 -5280 2630 -5210
rect 2590 -7137 2630 -6880
rect 2583 -7153 2637 -7137
rect 2583 -7187 2593 -7153
rect 2627 -7187 2637 -7153
rect 2583 -7203 2637 -7187
<< polycont >>
rect 2593 -7187 2627 -7153
<< locali >>
rect 2520 -6860 2530 -5184
rect 2520 -6880 2570 -6860
rect 2650 -5290 2700 -5190
rect 2650 -5310 2660 -5290
rect 2650 -6880 2700 -6860
rect 2590 -7153 2630 -7150
rect 2577 -7187 2593 -7153
rect 2627 -7187 2643 -7153
rect 2590 -7190 2630 -7187
<< viali >>
rect 2516 -5184 2604 -5096
rect 2530 -5310 2570 -5184
rect 2530 -6830 2570 -5310
rect 2660 -5310 2700 -5290
rect 2660 -6860 2690 -5310
rect 2690 -6860 2700 -5310
rect 2590 -7230 2630 -7190
<< metal1 >>
rect 2504 -4830 2510 -4730
rect 2610 -4830 2616 -4730
rect 2510 -5096 2520 -4830
rect 2600 -5096 2610 -4830
rect 2510 -5184 2516 -5096
rect 2604 -5184 2610 -5096
rect 2510 -6850 2520 -5184
rect 2600 -6850 2610 -5184
rect 2650 -5290 2730 -5190
rect 2650 -6860 2660 -5290
rect 2720 -6860 2730 -5290
rect 2650 -6880 2730 -6860
rect 2419 -6970 2770 -6920
rect 2440 -7020 2770 -6970
rect 2369 -7120 2770 -7020
rect 2584 -7184 2636 -7178
rect 2578 -7236 2584 -7184
rect 2636 -7236 2642 -7184
rect 2584 -7242 2636 -7236
<< via1 >>
rect 2510 -4830 2610 -4730
rect 2520 -5096 2600 -4830
rect 2520 -5184 2600 -5096
rect 2520 -6830 2530 -5184
rect 2530 -6830 2570 -5184
rect 2570 -6830 2600 -5184
rect 2520 -6850 2600 -6830
rect 2660 -6860 2700 -5290
rect 2700 -6860 2720 -5290
rect 2584 -7190 2636 -7184
rect 2584 -7230 2590 -7190
rect 2590 -7230 2630 -7190
rect 2630 -7230 2636 -7190
rect 2584 -7236 2636 -7230
<< metal2 >>
rect 939 -2920 969 -2860
rect 120 -2960 970 -2920
rect 1104 -2940 1144 -2860
rect 120 -3140 160 -2960
rect 1374 -3000 1404 -2860
rect 1539 -2940 1579 -2860
rect 940 -3040 1410 -3000
rect 1809 -3020 1839 -2860
rect 1974 -2940 2014 -2860
rect 359 -3060 419 -3051
rect 359 -3129 419 -3120
rect 29 -3180 160 -3140
rect 369 -3180 409 -3129
rect 940 -3140 980 -3040
rect 1480 -3060 1840 -3020
rect 1480 -3100 1520 -3060
rect 709 -3180 980 -3140
rect 1040 -3132 1130 -3110
rect 125 -3185 155 -3180
rect 1040 -3188 1062 -3132
rect 1118 -3188 1130 -3132
rect 1389 -3140 1520 -3100
rect 1690 -3113 1770 -3110
rect 1686 -3122 1770 -3113
rect 1389 -3180 1429 -3140
rect 1742 -3178 1770 -3122
rect 2244 -3140 2274 -2860
rect 2409 -2940 2449 -2860
rect 2399 -3040 2459 -3031
rect 2399 -3109 2459 -3100
rect 1686 -3187 1770 -3178
rect 2069 -3180 2274 -3140
rect 2409 -3180 2449 -3109
rect 2244 -3185 2274 -3180
rect 1040 -3210 1130 -3188
rect 1690 -3200 1770 -3187
rect 2510 -4730 2610 -4724
rect 2506 -4825 2510 -4735
rect 2610 -4825 2614 -4735
rect 2510 -6850 2520 -4830
rect 2600 -6850 2610 -4830
rect 2510 -6920 2610 -6850
rect 2650 -5240 2730 -5190
rect 2650 -6860 2660 -5240
rect 2720 -6860 2730 -5240
rect 2650 -6880 2730 -6860
rect 2580 -7180 2640 -7171
rect 2578 -7236 2580 -7184
rect 2640 -7236 2642 -7184
rect 2580 -7249 2640 -7240
<< via2 >>
rect 359 -3120 419 -3060
rect 1062 -3188 1118 -3132
rect 1686 -3178 1742 -3122
rect 2399 -3100 2459 -3040
rect 2515 -4825 2605 -4735
rect 2660 -5290 2720 -5240
rect 2660 -6070 2720 -5290
rect 2580 -7184 2640 -7180
rect 2580 -7236 2584 -7184
rect 2584 -7236 2636 -7184
rect 2636 -7236 2640 -7184
rect 2580 -7240 2640 -7236
<< metal3 >>
rect 2700 -2950 2800 -2930
rect 2380 -3035 2480 -3020
rect 350 -3055 550 -3040
rect 350 -3119 354 -3055
rect 424 -3119 550 -3055
rect 2380 -3099 2394 -3035
rect 2464 -3099 2480 -3035
rect 2380 -3100 2399 -3099
rect 2459 -3100 2480 -3099
rect 350 -3120 359 -3119
rect 419 -3120 550 -3119
rect 350 -3140 550 -3120
rect 1040 -3128 1160 -3110
rect 1040 -3192 1058 -3128
rect 1122 -3192 1160 -3128
rect 1040 -3210 1160 -3192
rect 1670 -3118 1790 -3110
rect 1670 -3182 1682 -3118
rect 1746 -3182 1790 -3118
rect 2380 -3130 2480 -3100
rect 1670 -3200 1790 -3182
rect 2700 -4720 2710 -2950
rect 2510 -4730 2710 -4720
rect 2510 -4731 2550 -4730
rect 2505 -4829 2511 -4731
rect 2510 -4830 2550 -4829
rect 2790 -4830 2800 -2950
rect 2510 -4840 2800 -4830
rect 2650 -5240 2730 -5190
rect 2650 -5520 2660 -5240
rect -770 -5920 2660 -5520
rect 2650 -6070 2660 -5920
rect 2720 -5520 2730 -5240
rect 2720 -5920 3480 -5520
rect 2720 -6070 2730 -5920
rect 2650 -6080 2730 -6070
rect 2550 -7180 2660 -7160
rect 2550 -7181 2580 -7180
rect 2640 -7181 2660 -7180
rect 2550 -7245 2575 -7181
rect 2645 -7245 2660 -7181
rect 2550 -7260 2660 -7245
<< via3 >>
rect 354 -3060 424 -3055
rect 354 -3119 359 -3060
rect 359 -3119 419 -3060
rect 419 -3119 424 -3060
rect 2394 -3040 2464 -3035
rect 2394 -3099 2399 -3040
rect 2399 -3099 2459 -3040
rect 2459 -3099 2464 -3040
rect 1058 -3132 1122 -3128
rect 1058 -3188 1062 -3132
rect 1062 -3188 1118 -3132
rect 1118 -3188 1122 -3132
rect 1058 -3192 1122 -3188
rect 1682 -3122 1746 -3118
rect 1682 -3178 1686 -3122
rect 1686 -3178 1742 -3122
rect 1742 -3178 1746 -3122
rect 1682 -3182 1746 -3178
rect 2710 -4730 2790 -2950
rect 2550 -4731 2790 -4730
rect 2511 -4735 2790 -4731
rect 2511 -4825 2515 -4735
rect 2515 -4825 2605 -4735
rect 2605 -4825 2790 -4735
rect 2511 -4829 2790 -4825
rect 2550 -4830 2790 -4829
rect 2575 -7240 2580 -7181
rect 2580 -7240 2640 -7181
rect 2640 -7240 2645 -7181
rect 2575 -7245 2645 -7240
<< metal4 >>
rect 353 -3055 425 -3054
rect 353 -3119 354 -3055
rect 424 -3060 425 -3055
rect 814 -3060 874 -2860
rect 1004 -2930 1064 -2860
rect 1249 -2880 1309 -2860
rect 424 -3119 874 -3060
rect 353 -3120 874 -3119
rect 1240 -2940 1309 -2880
rect 1439 -2940 1499 -2860
rect 1057 -3128 1123 -3127
rect 1057 -3192 1058 -3128
rect 1122 -3130 1123 -3128
rect 1240 -3130 1300 -2940
rect 1684 -3117 1744 -2860
rect 1874 -2940 1934 -2860
rect 2119 -3040 2179 -2860
rect 2309 -2940 2369 -2860
rect 2700 -2950 2800 -2860
rect 2393 -3035 2465 -3034
rect 2393 -3040 2394 -3035
rect 2119 -3099 2394 -3040
rect 2464 -3099 2465 -3035
rect 2119 -3100 2465 -3099
rect 1122 -3190 1300 -3130
rect 1681 -3118 1747 -3117
rect 1681 -3182 1682 -3118
rect 1746 -3182 1747 -3118
rect 1681 -3183 1747 -3182
rect 1122 -3192 1123 -3190
rect 1057 -3193 1123 -3192
rect 2700 -4720 2710 -2950
rect 2510 -4730 2710 -4720
rect 2510 -4731 2550 -4730
rect 2510 -4829 2511 -4731
rect 2510 -4830 2550 -4829
rect 2790 -4830 2800 -2950
rect 2510 -4840 2800 -4830
rect 2574 -7181 2646 -7180
rect 2574 -7245 2575 -7181
rect 2645 -7245 2646 -7181
rect 2574 -7246 2646 -7245
rect 2580 -7420 2640 -7246
use 8bit_sens  8bit_sens_0
timestamp 1662227450
transform 1 0 -251 0 1 -6480
box -110 -750 2810 3340
use pixel  pixel_0
timestamp 1662180122
transform 1 0 0 0 1 70
box -470 -3000 3090 570
<< labels >>
rlabel metal4 2341 -2908 2341 -2908 1 GRAYx1x
port 77 n
rlabel metal2 1989 -2907 1989 -2907 1 GRAYx2x
port 76 n
rlabel metal4 1903 -2922 1903 -2922 1 GRAYx3x
port 75 n
rlabel metal2 1553 -2891 1553 -2891 1 GRAYx4x
port 74 n
rlabel metal4 1470 -2911 1470 -2910 1 GRAYx5x
port 73 n
rlabel metal2 959 -2895 959 -2895 1 OUTx7x
port 72 n
rlabel metal4 841 -2921 841 -2921 1 OUTx6x
port 71 n
rlabel metal4 1031 -2900 1031 -2900 1 GRAYx7x
port 70 n
rlabel metal2 1119 -2906 1119 -2906 1 GRAYx6x
port 69 n
rlabel metal4 1283 -2898 1283 -2898 1 OUTx4x
port 68 n
rlabel metal2 1388 -2908 1388 -2908 1 OUTx5x
port 67 n
rlabel metal4 1716 -2898 1716 -2898 1 OUTx2x
port 64 n
rlabel metal2 1821 -2906 1821 -2906 1 OUTx3x
port 63 n
rlabel metal2 2256 -2915 2256 -2915 1 OUTx1x
port 59 n
rlabel metal2 2431 -2902 2431 -2902 1 GRAYx0x
port 57 n
rlabel metal4 2135 -2917 2135 -2917 1 OUTx0x
port 60 n
rlabel metal3 -730 -5710 -730 -5710 1 ARRAY_OUT
port 81 n
rlabel metal4 2600 -7340 2600 -7340 1 COL_SEL
port 82 n
<< end >>
