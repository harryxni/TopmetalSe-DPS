magic
tech sky130B
magscale 1 2
timestamp 1662181774
<< metal1 >>
rect -80 3120 4925 3270
rect 5075 3120 5081 3270
rect 3490 1590 5850 1650
rect 5910 1590 5916 1650
rect 3430 1355 4015 1505
rect 4165 1355 4171 1505
rect 3430 1025 3580 1355
rect 3430 875 3885 1025
rect 4035 875 4041 1025
rect 3430 480 3580 875
rect 90 330 420 480
rect 3085 330 3580 480
<< via1 >>
rect 4925 3120 5075 3270
rect 5850 1590 5910 1650
rect 4015 1355 4165 1505
rect 3885 875 4035 1025
<< metal2 >>
rect 4925 3270 5075 3276
rect 4916 3120 4925 3270
rect 5075 3120 5084 3270
rect 4925 3114 5075 3120
rect 5375 2098 5585 3645
rect 5375 2042 5452 2098
rect 5508 2042 5585 2098
rect 4015 1505 4165 1511
rect 4006 1355 4015 1505
rect 4165 1355 4174 1505
rect 4015 1349 4165 1355
rect 3885 1025 4035 1031
rect 3876 875 3885 1025
rect 4035 875 4044 1025
rect 3885 869 4035 875
rect 4379 738 4542 870
rect 4379 682 4432 738
rect 4488 682 4542 738
rect 4379 300 4542 682
rect 5375 -255 5585 2042
rect 5850 1650 5910 1659
rect 5850 1581 5910 1590
<< via2 >>
rect 4925 3120 5075 3270
rect 5452 2042 5508 2098
rect 4015 1355 4165 1505
rect 3885 875 4035 1025
rect 4432 682 4488 738
rect 5850 1590 5910 1650
<< metal3 >>
rect 4920 3270 4930 3275
rect 4920 3120 4925 3270
rect 4920 3115 4930 3120
rect 5080 3115 5086 3275
rect -80 2990 250 3050
rect -80 2790 60 2850
rect -80 2490 160 2550
rect 6608 2232 6672 2238
rect 3500 2170 6608 2230
rect 6608 2162 6672 2168
rect 5447 2100 5513 2103
rect 3470 2098 5513 2100
rect 3470 2042 5452 2098
rect 5508 2042 5513 2098
rect 3470 2040 5513 2042
rect 5447 2037 5513 2040
rect 6168 1932 6232 1938
rect 3500 1870 6168 1930
rect 6168 1862 6232 1868
rect 5820 1655 5930 1680
rect 5820 1591 5845 1655
rect 5915 1591 5930 1655
rect 5820 1590 5850 1591
rect 5910 1590 5930 1591
rect 5820 1560 5930 1590
rect 4010 1505 4020 1510
rect 4010 1355 4015 1505
rect 4010 1350 4020 1355
rect 4170 1350 4176 1510
rect 3880 1025 3890 1030
rect 3880 875 3885 1025
rect 3880 870 3890 875
rect 4040 870 4046 1030
rect 4427 740 4493 743
rect -80 680 80 740
rect 3470 738 4493 740
rect 3470 682 4432 738
rect 4488 682 4493 738
rect 3470 680 4493 682
rect 4427 677 4493 680
rect 4642 480 4648 482
rect 3500 420 4648 480
rect 4642 418 4648 420
rect 4712 418 4718 482
<< via3 >>
rect 4930 3270 5080 3275
rect 4930 3120 5075 3270
rect 5075 3120 5080 3270
rect 4930 3115 5080 3120
rect 6608 2168 6672 2232
rect 6168 1868 6232 1932
rect 5845 1650 5915 1655
rect 5845 1591 5850 1650
rect 5850 1591 5910 1650
rect 5910 1591 5915 1650
rect 4020 1505 4170 1510
rect 4020 1355 4165 1505
rect 4165 1355 4170 1505
rect 4020 1350 4170 1355
rect 3890 1025 4040 1030
rect 3890 875 4035 1025
rect 4035 875 4040 1025
rect 3890 870 4040 875
rect 4648 418 4712 482
<< metal4 >>
rect 3805 3160 4195 3640
rect 3835 3030 4185 3160
rect 4660 483 4720 3620
rect 4800 3490 5200 3650
rect 4800 3355 4855 3490
rect 5175 3370 5200 3490
rect 5175 3355 5210 3370
rect 4800 3035 4850 3355
rect 5180 3035 5210 3355
rect 4800 2820 4855 3035
rect 5175 3030 5210 3035
rect 5175 2820 5200 3030
rect 5850 1656 5910 3640
rect 6170 1933 6230 3640
rect 6460 3455 6840 3560
rect 6460 2360 6500 3455
rect 6460 2040 6480 2360
rect 6167 1932 6233 1933
rect 6167 1868 6168 1932
rect 6232 1868 6233 1932
rect 6167 1867 6233 1868
rect 5844 1655 5916 1656
rect 5844 1591 5845 1655
rect 5915 1591 5916 1655
rect 5844 1590 5916 1591
rect 4647 482 4720 483
rect 4647 418 4648 482
rect 4712 418 4720 482
rect 4647 417 4720 418
rect 4660 -50 4720 417
rect 4830 110 5190 290
rect 5850 -220 5910 1590
rect 6170 -270 6230 1867
rect 6460 570 6500 2040
rect 6810 570 6840 3455
rect 6460 -310 6840 570
<< via4 >>
rect 3855 1590 4175 3030
rect 3855 1510 4255 1590
rect 3855 1350 4020 1510
rect 4020 1350 4170 1510
rect 4170 1350 4255 1510
rect 3855 1270 4255 1350
rect 3855 1110 4175 1270
rect 3805 1030 4175 1110
rect 3805 870 3890 1030
rect 3890 870 4040 1030
rect 4040 870 4175 1030
rect 3805 790 4175 870
rect 3855 170 4175 790
rect 4855 3355 5175 3490
rect 4850 3275 5180 3355
rect 4850 3115 4930 3275
rect 4930 3115 5080 3275
rect 5080 3115 5180 3275
rect 4850 3035 5180 3115
rect 4855 650 5175 3035
rect 6500 2360 6810 3455
rect 6480 2232 6810 2360
rect 6480 2168 6608 2232
rect 6608 2168 6672 2232
rect 6672 2168 6810 2232
rect 6480 2040 6810 2168
rect 6500 570 6810 2040
<< metal5 >>
rect 3805 3320 4195 3640
rect 4800 3490 5200 3650
rect 4800 3355 4855 3490
rect 5175 3379 5200 3490
rect 6460 3455 6840 3630
rect 5175 3355 5213 3379
rect 3805 3030 4205 3320
rect 3805 1134 3855 3030
rect 4175 1614 4205 3030
rect 4800 3035 4850 3355
rect 5180 3035 5213 3355
rect 4800 2820 4855 3035
rect 4175 1590 4279 1614
rect 4255 1270 4279 1590
rect 3781 1110 3855 1134
rect 4175 1246 4279 1270
rect 3781 790 3805 1110
rect 3781 766 3855 790
rect 3805 170 3855 766
rect 4175 170 4205 1246
rect 3805 -120 4205 170
rect 4805 650 4855 2820
rect 5175 3011 5213 3035
rect 5175 650 5205 3011
rect 6460 2384 6500 3455
rect 6456 2360 6500 2384
rect 6456 2040 6480 2360
rect 6456 2016 6500 2040
rect 4805 -120 5205 650
rect 6460 570 6500 2016
rect 6810 570 6840 3455
rect 6460 -310 6840 570
use pixel  pixel_0
timestamp 1662180122
transform 1 0 470 0 1 3000
box -470 -3000 3090 570
<< end >>
