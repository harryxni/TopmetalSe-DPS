magic
tech sky130B
magscale 1 2
timestamp 1662068818
<< nwell >>
rect 1920 290 2800 300
rect -200 -60 2800 290
rect -200 -370 1920 -60
rect 960 -1180 2385 -750
<< pwell >>
rect 2424 -164 2616 -154
rect 2364 -324 2616 -164
rect 464 -454 716 -414
rect -166 -806 716 -454
rect 2174 -706 2626 -324
rect -56 -1236 526 -806
rect -56 -2374 236 -1236
rect 974 -1314 1196 -1224
rect 1594 -1304 1816 -1224
rect 2134 -1304 2366 -1224
rect 1594 -1314 2366 -1304
rect 974 -1476 2366 -1314
rect 1304 -1716 1456 -1476
rect 1844 -1696 2096 -1476
rect -56 -2666 416 -2374
<< nmos >>
rect 1330 -1620 1420 -1420
rect 2230 -1450 2260 -1250
<< pmos >>
rect 2220 -1110 2260 -910
<< pmoslvt >>
rect -50 10 350 210
rect 420 10 820 210
rect 1060 10 1460 210
rect 1530 10 1930 210
rect 2130 -20 2330 180
rect 2430 -20 2630 180
rect 120 -320 1720 -236
rect 1070 -1060 1270 -860
rect 1520 -1060 1720 -860
rect 1930 -1060 2020 -860
<< nmoslvt >>
rect 2390 -280 2590 -250
rect -140 -710 60 -550
rect 120 -710 320 -550
rect 490 -710 690 -510
rect 2200 -580 2600 -380
rect 20 -2250 50 -850
rect 130 -2250 160 -850
rect 300 -1130 500 -890
rect 1070 -1450 1100 -1250
rect 1690 -1450 1720 -1250
rect 1870 -1600 2070 -1400
rect 40 -2640 240 -2400
<< ndiff >>
rect 2450 -190 2590 -180
rect 2390 -193 2590 -190
rect 2390 -227 2503 -193
rect 2537 -227 2590 -193
rect 2390 -250 2590 -227
rect 2390 -350 2590 -280
rect 2200 -380 2600 -350
rect 490 -453 690 -440
rect -140 -493 60 -480
rect -140 -527 -91 -493
rect -57 -527 -23 -493
rect 11 -527 60 -493
rect -140 -550 60 -527
rect 120 -493 320 -480
rect 120 -527 169 -493
rect 203 -527 237 -493
rect 271 -527 320 -493
rect 490 -487 539 -453
rect 573 -487 607 -453
rect 641 -487 690 -453
rect 490 -510 690 -487
rect 120 -550 320 -527
rect 2200 -623 2600 -580
rect 2200 -657 2247 -623
rect 2281 -657 2315 -623
rect 2349 -657 2383 -623
rect 2417 -657 2451 -623
rect 2485 -657 2519 -623
rect 2553 -657 2600 -623
rect 2200 -680 2600 -657
rect -140 -780 60 -710
rect 120 -780 320 -710
rect 490 -730 690 -710
rect 460 -733 690 -730
rect 460 -767 539 -733
rect 573 -767 607 -733
rect 641 -767 690 -733
rect 460 -780 690 -767
rect -30 -850 0 -780
rect 180 -850 210 -780
rect 460 -840 500 -780
rect -30 -2250 20 -850
rect 50 -911 130 -850
rect 50 -945 73 -911
rect 107 -945 130 -911
rect 50 -979 130 -945
rect 50 -1013 73 -979
rect 107 -1013 130 -979
rect 50 -1047 130 -1013
rect 50 -1081 73 -1047
rect 107 -1081 130 -1047
rect 50 -1115 130 -1081
rect 50 -1149 73 -1115
rect 107 -1149 130 -1115
rect 50 -1183 130 -1149
rect 50 -1217 73 -1183
rect 107 -1217 130 -1183
rect 50 -1251 130 -1217
rect 50 -1285 73 -1251
rect 107 -1285 130 -1251
rect 50 -1319 130 -1285
rect 50 -1353 73 -1319
rect 107 -1353 130 -1319
rect 50 -1387 130 -1353
rect 50 -1421 73 -1387
rect 107 -1421 130 -1387
rect 50 -1455 130 -1421
rect 50 -1489 73 -1455
rect 107 -1489 130 -1455
rect 50 -1523 130 -1489
rect 50 -1557 73 -1523
rect 107 -1557 130 -1523
rect 50 -1591 130 -1557
rect 50 -1625 73 -1591
rect 107 -1625 130 -1591
rect 50 -1659 130 -1625
rect 50 -1693 73 -1659
rect 107 -1693 130 -1659
rect 50 -1727 130 -1693
rect 50 -1761 73 -1727
rect 107 -1761 130 -1727
rect 50 -1795 130 -1761
rect 50 -1829 73 -1795
rect 107 -1829 130 -1795
rect 50 -1863 130 -1829
rect 50 -1897 73 -1863
rect 107 -1897 130 -1863
rect 50 -1931 130 -1897
rect 50 -1965 73 -1931
rect 107 -1965 130 -1931
rect 50 -1999 130 -1965
rect 50 -2033 73 -1999
rect 107 -2033 130 -1999
rect 50 -2067 130 -2033
rect 50 -2101 73 -2067
rect 107 -2101 130 -2067
rect 50 -2135 130 -2101
rect 50 -2169 73 -2135
rect 107 -2169 130 -2135
rect 50 -2250 130 -2169
rect 160 -2250 210 -850
rect 300 -890 500 -840
rect 300 -1158 500 -1130
rect 300 -1192 349 -1158
rect 383 -1192 417 -1158
rect 451 -1192 500 -1158
rect 300 -1210 500 -1192
rect 1000 -1299 1070 -1250
rect 1000 -1333 1013 -1299
rect 1047 -1333 1070 -1299
rect 1000 -1367 1070 -1333
rect 1000 -1401 1013 -1367
rect 1047 -1401 1070 -1367
rect 1000 -1450 1070 -1401
rect 1100 -1299 1170 -1250
rect 1100 -1333 1123 -1299
rect 1157 -1333 1170 -1299
rect 1100 -1367 1170 -1333
rect 1620 -1299 1690 -1250
rect 1620 -1333 1633 -1299
rect 1667 -1333 1690 -1299
rect 1100 -1401 1123 -1367
rect 1157 -1401 1170 -1367
rect 1100 -1450 1170 -1401
rect 1330 -1358 1420 -1340
rect 1330 -1392 1358 -1358
rect 1392 -1392 1420 -1358
rect 1330 -1420 1420 -1392
rect 1620 -1367 1690 -1333
rect 1620 -1401 1633 -1367
rect 1667 -1401 1690 -1367
rect 1620 -1450 1690 -1401
rect 1720 -1299 1790 -1250
rect 1720 -1333 1743 -1299
rect 1777 -1333 1790 -1299
rect 2160 -1299 2230 -1250
rect 1720 -1367 1790 -1333
rect 1720 -1401 1743 -1367
rect 1777 -1401 1790 -1367
rect 1870 -1343 2070 -1330
rect 1870 -1377 1919 -1343
rect 1953 -1377 1987 -1343
rect 2021 -1377 2070 -1343
rect 1870 -1400 2070 -1377
rect 2160 -1333 2173 -1299
rect 2207 -1333 2230 -1299
rect 2160 -1367 2230 -1333
rect 1720 -1450 1790 -1401
rect 2160 -1401 2173 -1367
rect 2207 -1401 2230 -1367
rect 2160 -1450 2230 -1401
rect 2260 -1299 2340 -1250
rect 2260 -1333 2288 -1299
rect 2322 -1333 2340 -1299
rect 2260 -1367 2340 -1333
rect 2260 -1401 2288 -1367
rect 2322 -1401 2340 -1367
rect 2260 -1450 2340 -1401
rect 1330 -1640 1420 -1620
rect 1870 -1623 2070 -1600
rect 1330 -1643 1430 -1640
rect 1330 -1677 1373 -1643
rect 1407 -1677 1430 -1643
rect 1870 -1657 1924 -1623
rect 1958 -1657 1992 -1623
rect 2026 -1657 2070 -1623
rect 1870 -1670 2070 -1657
rect 1330 -1690 1430 -1677
rect -30 -2430 40 -2400
rect -30 -2464 -17 -2430
rect 17 -2464 40 -2430
rect -30 -2498 40 -2464
rect -30 -2532 -17 -2498
rect 17 -2532 40 -2498
rect -30 -2566 40 -2532
rect -30 -2600 -17 -2566
rect 17 -2600 40 -2566
rect -30 -2640 40 -2600
rect 240 -2430 310 -2400
rect 240 -2464 263 -2430
rect 297 -2464 310 -2430
rect 240 -2498 310 -2464
rect 240 -2532 263 -2498
rect 297 -2532 310 -2498
rect 240 -2566 310 -2532
rect 240 -2600 263 -2566
rect 297 -2600 310 -2566
rect 240 -2640 310 -2600
<< pdiff >>
rect -120 141 -50 210
rect -120 107 -107 141
rect -73 107 -50 141
rect -120 73 -50 107
rect -120 39 -107 73
rect -73 39 -50 73
rect -120 10 -50 39
rect 350 134 420 210
rect 350 100 370 134
rect 404 100 420 134
rect 350 54 420 100
rect 350 20 370 54
rect 404 20 420 54
rect 350 10 420 20
rect 820 161 890 210
rect 990 161 1060 210
rect 820 127 843 161
rect 877 127 890 161
rect 990 127 1003 161
rect 1037 127 1060 161
rect 820 93 890 127
rect 990 93 1060 127
rect 820 59 843 93
rect 877 59 890 93
rect 990 59 1003 93
rect 1037 59 1060 93
rect 820 10 890 59
rect 990 10 1060 59
rect 1460 10 1530 210
rect 1930 134 2000 210
rect 1930 100 1950 134
rect 1984 100 2000 134
rect 1930 54 2000 100
rect 1930 20 1950 54
rect 1984 20 2000 54
rect 1930 10 2000 20
rect 2060 129 2130 180
rect 2060 95 2076 129
rect 2110 95 2130 129
rect 2060 61 2130 95
rect 2060 27 2076 61
rect 2110 27 2130 61
rect 2060 -20 2130 27
rect 2330 121 2430 180
rect 2330 87 2363 121
rect 2397 87 2430 121
rect 2330 53 2430 87
rect 2330 19 2363 53
rect 2397 19 2430 53
rect 2330 -20 2430 19
rect 2630 131 2700 180
rect 2630 97 2653 131
rect 2687 97 2700 131
rect 2630 63 2700 97
rect 2630 29 2653 63
rect 2687 29 2700 63
rect 2630 -20 2700 29
rect -10 -268 120 -236
rect -10 -302 33 -268
rect 67 -302 120 -268
rect -10 -320 120 -302
rect 1720 -255 1860 -236
rect 1720 -289 1768 -255
rect 1802 -289 1860 -255
rect 1720 -320 1860 -289
rect 1000 -909 1070 -860
rect 1000 -943 1013 -909
rect 1047 -943 1070 -909
rect 1000 -977 1070 -943
rect 1000 -1011 1013 -977
rect 1047 -1011 1070 -977
rect 1000 -1060 1070 -1011
rect 1270 -909 1350 -860
rect 1450 -909 1520 -860
rect 1270 -943 1293 -909
rect 1327 -943 1350 -909
rect 1450 -943 1471 -909
rect 1505 -943 1520 -909
rect 1270 -977 1350 -943
rect 1450 -977 1520 -943
rect 1270 -1011 1293 -977
rect 1327 -1011 1350 -977
rect 1450 -1011 1471 -977
rect 1505 -1011 1520 -977
rect 1270 -1060 1350 -1011
rect 1450 -1060 1520 -1011
rect 1720 -909 1790 -860
rect 1720 -943 1743 -909
rect 1777 -943 1790 -909
rect 1720 -977 1790 -943
rect 1720 -1011 1743 -977
rect 1777 -1011 1790 -977
rect 1720 -1060 1790 -1011
rect 1860 -909 1930 -860
rect 1860 -943 1873 -909
rect 1907 -943 1930 -909
rect 1860 -977 1930 -943
rect 1860 -1011 1873 -977
rect 1907 -1011 1930 -977
rect 1860 -1060 1930 -1011
rect 2020 -909 2090 -860
rect 2020 -943 2043 -909
rect 2077 -943 2090 -909
rect 2020 -977 2090 -943
rect 2020 -1011 2043 -977
rect 2077 -1011 2090 -977
rect 2020 -1060 2090 -1011
rect 2150 -959 2220 -910
rect 2150 -993 2166 -959
rect 2200 -993 2220 -959
rect 2150 -1027 2220 -993
rect 2150 -1061 2166 -1027
rect 2200 -1061 2220 -1027
rect 2150 -1110 2220 -1061
rect 2260 -959 2330 -910
rect 2260 -993 2283 -959
rect 2317 -993 2330 -959
rect 2260 -1027 2330 -993
rect 2260 -1061 2283 -1027
rect 2317 -1061 2330 -1027
rect 2260 -1110 2330 -1061
<< ndiffc >>
rect 2503 -227 2537 -193
rect -91 -527 -57 -493
rect -23 -527 11 -493
rect 169 -527 203 -493
rect 237 -527 271 -493
rect 539 -487 573 -453
rect 607 -487 641 -453
rect 2247 -657 2281 -623
rect 2315 -657 2349 -623
rect 2383 -657 2417 -623
rect 2451 -657 2485 -623
rect 2519 -657 2553 -623
rect 539 -767 573 -733
rect 607 -767 641 -733
rect 73 -945 107 -911
rect 73 -1013 107 -979
rect 73 -1081 107 -1047
rect 73 -1149 107 -1115
rect 73 -1217 107 -1183
rect 73 -1285 107 -1251
rect 73 -1353 107 -1319
rect 73 -1421 107 -1387
rect 73 -1489 107 -1455
rect 73 -1557 107 -1523
rect 73 -1625 107 -1591
rect 73 -1693 107 -1659
rect 73 -1761 107 -1727
rect 73 -1829 107 -1795
rect 73 -1897 107 -1863
rect 73 -1965 107 -1931
rect 73 -2033 107 -1999
rect 73 -2101 107 -2067
rect 73 -2169 107 -2135
rect 349 -1192 383 -1158
rect 417 -1192 451 -1158
rect 1013 -1333 1047 -1299
rect 1013 -1401 1047 -1367
rect 1123 -1333 1157 -1299
rect 1633 -1333 1667 -1299
rect 1123 -1401 1157 -1367
rect 1358 -1392 1392 -1358
rect 1633 -1401 1667 -1367
rect 1743 -1333 1777 -1299
rect 1743 -1401 1777 -1367
rect 1919 -1377 1953 -1343
rect 1987 -1377 2021 -1343
rect 2173 -1333 2207 -1299
rect 2173 -1401 2207 -1367
rect 2288 -1333 2322 -1299
rect 2288 -1401 2322 -1367
rect 1373 -1677 1407 -1643
rect 1924 -1657 1958 -1623
rect 1992 -1657 2026 -1623
rect -17 -2464 17 -2430
rect -17 -2532 17 -2498
rect -17 -2600 17 -2566
rect 263 -2464 297 -2430
rect 263 -2532 297 -2498
rect 263 -2600 297 -2566
<< pdiffc >>
rect -107 107 -73 141
rect -107 39 -73 73
rect 370 100 404 134
rect 370 20 404 54
rect 843 127 877 161
rect 1003 127 1037 161
rect 843 59 877 93
rect 1003 59 1037 93
rect 1950 100 1984 134
rect 1950 20 1984 54
rect 2076 95 2110 129
rect 2076 27 2110 61
rect 2363 87 2397 121
rect 2363 19 2397 53
rect 2653 97 2687 131
rect 2653 29 2687 63
rect 33 -302 67 -268
rect 1768 -289 1802 -255
rect 1013 -943 1047 -909
rect 1013 -1011 1047 -977
rect 1293 -943 1327 -909
rect 1471 -943 1505 -909
rect 1293 -1011 1327 -977
rect 1471 -1011 1505 -977
rect 1743 -943 1777 -909
rect 1743 -1011 1777 -977
rect 1873 -943 1907 -909
rect 1873 -1011 1907 -977
rect 2043 -943 2077 -909
rect 2043 -1011 2077 -977
rect 2166 -993 2200 -959
rect 2166 -1061 2200 -1027
rect 2283 -993 2317 -959
rect 2283 -1061 2317 -1027
<< psubdiff >>
rect 310 -2435 390 -2400
rect 310 -2469 343 -2435
rect 377 -2469 390 -2435
rect 310 -2503 390 -2469
rect 310 -2537 343 -2503
rect 377 -2537 390 -2503
rect 310 -2571 390 -2537
rect 310 -2605 343 -2571
rect 377 -2605 390 -2571
rect 310 -2640 390 -2605
<< nsubdiff >>
rect 890 161 990 210
rect 890 127 923 161
rect 957 127 990 161
rect 890 93 990 127
rect 890 59 923 93
rect 957 59 990 93
rect 890 10 990 59
rect 1350 -909 1450 -860
rect 1350 -943 1383 -909
rect 1417 -943 1450 -909
rect 1350 -977 1450 -943
rect 1350 -1011 1383 -977
rect 1417 -1011 1450 -977
rect 1350 -1060 1450 -1011
<< psubdiffcont >>
rect 343 -2469 377 -2435
rect 343 -2537 377 -2503
rect 343 -2605 377 -2571
<< nsubdiffcont >>
rect 923 127 957 161
rect 923 59 957 93
rect 1383 -943 1417 -909
rect 1383 -1011 1417 -977
<< poly >>
rect -50 210 350 240
rect 420 210 820 240
rect 1060 210 1460 240
rect 1530 210 1930 240
rect 2130 180 2330 210
rect 2430 180 2630 210
rect -50 -20 350 10
rect 420 -20 820 10
rect 1060 -20 1460 10
rect 1530 -20 1930 10
rect -10 -53 70 -20
rect -10 -87 8 -53
rect 42 -87 70 -53
rect -10 -110 70 -87
rect 480 -43 560 -20
rect 480 -77 503 -43
rect 537 -77 560 -43
rect 770 -50 1110 -20
rect 1530 -50 1600 -20
rect 2130 -50 2330 -20
rect 2430 -50 2630 -20
rect 480 -90 560 -77
rect 1530 -63 1590 -50
rect 1530 -97 1543 -63
rect 1577 -97 1590 -63
rect 1530 -116 1590 -97
rect 2130 -98 2210 -50
rect 2430 -73 2520 -50
rect 2430 -80 2463 -73
rect 1230 -143 1340 -130
rect 1230 -177 1273 -143
rect 1307 -177 1340 -143
rect 2130 -132 2153 -98
rect 2187 -132 2210 -98
rect 2440 -107 2463 -80
rect 2497 -107 2520 -73
rect 2440 -120 2520 -107
rect 2130 -160 2210 -132
rect 1230 -208 1340 -177
rect 120 -236 1720 -208
rect 2287 -248 2353 -238
rect 2287 -282 2303 -248
rect 2337 -250 2353 -248
rect 2337 -280 2390 -250
rect 2590 -280 2620 -250
rect 2337 -282 2353 -280
rect 2287 -292 2353 -282
rect 120 -350 1720 -320
rect -200 -710 -140 -550
rect 60 -710 120 -550
rect 320 -710 350 -550
rect 400 -559 490 -510
rect 400 -593 413 -559
rect 447 -593 490 -559
rect 400 -627 490 -593
rect 400 -661 413 -627
rect 447 -661 490 -627
rect 400 -710 490 -661
rect 690 -710 720 -510
rect 2170 -580 2200 -380
rect 2600 -398 2720 -380
rect 2600 -432 2658 -398
rect 2692 -432 2720 -398
rect 2600 -460 2720 -432
rect 2600 -580 2630 -460
rect -200 -850 -170 -710
rect 20 -850 50 -820
rect 130 -850 160 -820
rect -200 -893 -130 -850
rect -200 -903 -97 -893
rect -200 -937 -147 -903
rect -113 -937 -97 -903
rect -200 -947 -97 -937
rect -200 -950 -130 -947
rect -150 -2268 -60 -2240
rect 1070 -860 1270 -830
rect 1520 -860 1720 -830
rect 1930 -860 2020 -830
rect 270 -1130 300 -890
rect 500 -1070 530 -890
rect 2220 -910 2260 -880
rect 500 -1083 630 -1070
rect 500 -1117 558 -1083
rect 592 -1117 630 -1083
rect 500 -1130 630 -1117
rect 1070 -1090 1270 -1060
rect 1520 -1090 1720 -1060
rect 1930 -1090 2020 -1060
rect 1070 -1123 1150 -1090
rect 1070 -1157 1093 -1123
rect 1127 -1157 1150 -1123
rect 1235 -1130 1550 -1090
rect 1930 -1107 1980 -1090
rect 1918 -1123 1980 -1107
rect 1680 -1143 1720 -1140
rect 1070 -1170 1150 -1157
rect 1617 -1153 1720 -1143
rect 1617 -1187 1633 -1153
rect 1667 -1187 1720 -1153
rect 1918 -1157 1928 -1123
rect 1962 -1157 1980 -1123
rect 2220 -1150 2260 -1110
rect 1918 -1170 1980 -1157
rect 1918 -1173 1972 -1170
rect 1617 -1197 1720 -1187
rect 1680 -1200 1720 -1197
rect 1070 -1250 1100 -1220
rect 1690 -1250 1720 -1200
rect 2027 -1193 2093 -1183
rect 2027 -1227 2043 -1193
rect 2077 -1195 2093 -1193
rect 2230 -1195 2260 -1150
rect 2077 -1225 2260 -1195
rect 2077 -1227 2093 -1225
rect 2027 -1237 2093 -1227
rect 2230 -1250 2260 -1225
rect 1250 -1440 1330 -1420
rect 1070 -1497 1100 -1450
rect 1240 -1489 1330 -1440
rect 1058 -1513 1112 -1497
rect 1058 -1547 1068 -1513
rect 1102 -1547 1112 -1513
rect 1058 -1563 1112 -1547
rect 1240 -1523 1253 -1489
rect 1287 -1523 1330 -1489
rect 1240 -1557 1330 -1523
rect 1240 -1591 1253 -1557
rect 1287 -1591 1330 -1557
rect 1240 -1620 1330 -1591
rect 1420 -1620 1460 -1420
rect 1690 -1480 1720 -1450
rect 1840 -1520 1870 -1400
rect 1770 -1548 1870 -1520
rect 1770 -1582 1793 -1548
rect 1827 -1582 1870 -1548
rect 1770 -1600 1870 -1582
rect 2070 -1600 2100 -1400
rect 2230 -1500 2260 -1450
rect 1770 -1610 1840 -1600
rect 230 -2193 330 -2160
rect 230 -2227 263 -2193
rect 297 -2227 330 -2193
rect -150 -2302 -122 -2268
rect -88 -2270 -60 -2268
rect 20 -2270 50 -2250
rect -88 -2300 50 -2270
rect 130 -2270 160 -2250
rect 230 -2270 330 -2227
rect 130 -2300 330 -2270
rect -88 -2302 -60 -2300
rect -150 -2330 -60 -2302
rect 453 -2348 507 -2332
rect 453 -2350 463 -2348
rect 180 -2370 463 -2350
rect 40 -2380 463 -2370
rect 40 -2400 240 -2380
rect 453 -2382 463 -2380
rect 497 -2382 507 -2348
rect 453 -2398 507 -2382
rect 40 -2670 240 -2640
<< polycont >>
rect 8 -87 42 -53
rect 503 -77 537 -43
rect 1543 -97 1577 -63
rect 1273 -177 1307 -143
rect 2153 -132 2187 -98
rect 2463 -107 2497 -73
rect 2303 -282 2337 -248
rect 413 -593 447 -559
rect 413 -661 447 -627
rect 2658 -432 2692 -398
rect -147 -937 -113 -903
rect 558 -1117 592 -1083
rect 1093 -1157 1127 -1123
rect 1633 -1187 1667 -1153
rect 1928 -1157 1962 -1123
rect 2043 -1227 2077 -1193
rect 1068 -1547 1102 -1513
rect 1253 -1523 1287 -1489
rect 1253 -1591 1287 -1557
rect 1793 -1582 1827 -1548
rect 263 -2227 297 -2193
rect -122 -2302 -88 -2268
rect 463 -2382 497 -2348
<< locali >>
rect 890 252 990 270
rect 2650 260 2690 270
rect 890 218 923 252
rect 957 218 990 252
rect 2630 257 2710 260
rect 2630 223 2653 257
rect 2687 223 2710 257
rect 2630 220 2710 223
rect 890 210 990 218
rect -120 141 -70 170
rect -120 107 -107 141
rect -73 107 -70 141
rect -120 73 -70 107
rect -120 39 -107 73
rect -73 39 -70 73
rect -120 -50 -70 39
rect 370 134 410 210
rect 404 100 410 134
rect 370 54 410 100
rect 404 20 410 54
rect -10 -50 70 -10
rect -120 -53 70 -50
rect -120 -87 8 -53
rect 42 -87 70 -53
rect 370 -30 410 20
rect 820 161 1060 210
rect 820 127 843 161
rect 877 127 923 161
rect 957 127 1003 161
rect 1037 127 1060 161
rect 820 93 1060 127
rect 820 59 843 93
rect 877 59 923 93
rect 957 59 1003 93
rect 1037 59 1060 93
rect 820 10 1060 59
rect 1950 134 1990 210
rect 1984 100 1990 134
rect 1950 54 1990 100
rect 1984 20 1990 54
rect 480 -30 560 -10
rect 370 -43 560 -30
rect 370 -70 503 -43
rect -120 -100 70 -87
rect 480 -77 503 -70
rect 537 -77 560 -43
rect 480 -90 560 -77
rect 1084 -60 1590 -50
rect 1084 -63 1596 -60
rect 1084 -90 1543 -63
rect -120 -400 -70 -100
rect -10 -110 70 -100
rect 30 -150 70 -110
rect 1084 -150 1124 -90
rect 1520 -97 1543 -90
rect 1577 -97 1596 -63
rect 1520 -100 1596 -97
rect 1520 -120 1590 -100
rect 1520 -121 1589 -120
rect 30 -190 1124 -150
rect 1220 -143 1350 -130
rect 1950 -140 1990 20
rect 1220 -160 1273 -143
rect 1180 -163 1273 -160
rect 1180 -197 1183 -163
rect 1217 -177 1273 -163
rect 1307 -177 1350 -143
rect 1217 -197 1350 -177
rect 1180 -200 1350 -197
rect 1630 -180 1990 -140
rect 2030 129 2110 180
rect 2030 95 2076 129
rect 2030 61 2110 95
rect 2030 27 2076 61
rect 2030 -20 2110 27
rect 2350 121 2410 170
rect 2350 87 2363 121
rect 2397 87 2410 121
rect 2350 53 2410 87
rect 2350 19 2363 53
rect 2397 19 2410 53
rect 2030 -163 2080 -20
rect 2120 -98 2220 -80
rect 2120 -132 2153 -98
rect 2187 -132 2220 -98
rect 2350 -100 2410 19
rect 2650 131 2690 220
rect 2650 97 2653 131
rect 2687 97 2690 131
rect 2650 63 2690 97
rect 2650 29 2653 63
rect 2687 29 2690 63
rect 2120 -160 2220 -132
rect 2300 -140 2410 -100
rect 2450 -73 2540 -50
rect 2450 -107 2463 -73
rect 2497 -78 2540 -73
rect 2450 -112 2473 -107
rect 2507 -112 2540 -78
rect 2450 -130 2540 -112
rect -10 -268 110 -250
rect -10 -302 33 -268
rect 67 -302 110 -268
rect 1630 -270 1670 -180
rect 2030 -197 2038 -163
rect 2072 -197 2080 -163
rect 2030 -220 2080 -197
rect -10 -320 110 -302
rect 280 -310 1670 -270
rect 1740 -255 1830 -236
rect 1740 -289 1768 -255
rect 1802 -260 1830 -255
rect 2130 -260 2210 -160
rect 1802 -289 2210 -260
rect -10 -383 60 -320
rect -120 -441 -71 -400
rect -10 -417 8 -383
rect 42 -417 60 -383
rect -10 -435 60 -417
rect 280 -430 320 -310
rect 1740 -320 2210 -289
rect 2300 -248 2340 -140
rect 2650 -180 2690 29
rect 2450 -193 2690 -180
rect 2450 -227 2503 -193
rect 2537 -227 2690 -193
rect 2450 -230 2690 -227
rect 2300 -282 2303 -248
rect 2337 -282 2340 -248
rect 2300 -300 2340 -282
rect 1740 -370 1790 -320
rect 500 -393 680 -390
rect 500 -427 537 -393
rect 571 -427 609 -393
rect 643 -427 680 -393
rect -120 -460 -70 -441
rect -140 -480 -70 -460
rect 280 -470 450 -430
rect 280 -480 320 -470
rect -140 -493 60 -480
rect -140 -527 -91 -493
rect -57 -527 -23 -493
rect 11 -527 60 -493
rect -140 -540 60 -527
rect 120 -493 320 -480
rect 120 -527 169 -493
rect 203 -527 237 -493
rect 271 -527 320 -493
rect 120 -540 320 -527
rect 400 -510 450 -470
rect 500 -453 680 -427
rect 500 -487 539 -453
rect 573 -487 607 -453
rect 641 -487 680 -453
rect 500 -510 680 -487
rect 740 -410 1790 -370
rect 2640 -388 2710 -360
rect 400 -559 460 -510
rect 400 -593 413 -559
rect 447 -593 460 -559
rect 400 -627 460 -593
rect 400 -661 413 -627
rect 447 -661 460 -627
rect 400 -710 460 -661
rect 490 -733 690 -730
rect 490 -743 539 -733
rect 573 -743 607 -733
rect 490 -777 517 -743
rect 573 -767 589 -743
rect 641 -750 690 -733
rect 740 -750 780 -410
rect 2640 -432 2658 -388
rect 2692 -432 2710 -388
rect 2640 -470 2710 -432
rect 2200 -620 2600 -600
rect 2200 -623 2690 -620
rect 2200 -657 2247 -623
rect 2281 -657 2315 -623
rect 2349 -657 2383 -623
rect 2417 -657 2451 -623
rect 2485 -657 2519 -623
rect 2553 -633 2690 -623
rect 2553 -657 2643 -633
rect 2200 -667 2643 -657
rect 2677 -667 2690 -633
rect 2200 -680 2690 -667
rect 2200 -690 2600 -680
rect 1350 -740 1450 -730
rect 641 -767 780 -750
rect 551 -777 589 -767
rect 623 -777 780 -767
rect 490 -790 780 -777
rect 1100 -758 2270 -740
rect 1100 -792 1179 -758
rect 1213 -792 1251 -758
rect 1285 -792 1323 -758
rect 1357 -792 1395 -758
rect 1429 -792 1467 -758
rect 1501 -792 1539 -758
rect 1573 -792 1611 -758
rect 1645 -792 1683 -758
rect 1717 -792 1755 -758
rect 1789 -792 1827 -758
rect 1861 -792 1899 -758
rect 1933 -792 1971 -758
rect 2005 -792 2043 -758
rect 2077 -792 2115 -758
rect 2149 -792 2187 -758
rect 2221 -792 2270 -758
rect 1100 -810 2270 -792
rect -147 -903 -113 -887
rect -147 -953 -113 -937
rect 60 -911 120 -850
rect 1350 -860 1450 -810
rect 60 -945 73 -911
rect 107 -945 120 -911
rect 60 -979 120 -945
rect 1000 -909 1050 -860
rect 1000 -943 1013 -909
rect 1047 -943 1050 -909
rect 60 -1013 73 -979
rect 107 -1013 120 -979
rect 60 -1047 120 -1013
rect 60 -1081 73 -1047
rect 107 -1081 120 -1047
rect 590 -963 630 -960
rect 590 -997 593 -963
rect 627 -997 630 -963
rect 590 -1070 630 -997
rect 1000 -977 1050 -943
rect 1000 -1011 1013 -977
rect 1047 -1011 1050 -977
rect 60 -1115 120 -1081
rect 60 -1149 73 -1115
rect 107 -1149 120 -1115
rect 530 -1083 630 -1070
rect 530 -1117 558 -1083
rect 592 -1117 630 -1083
rect 530 -1130 630 -1117
rect 800 -1033 870 -1015
rect 800 -1067 818 -1033
rect 852 -1067 870 -1033
rect 60 -1183 120 -1149
rect 60 -1217 73 -1183
rect 107 -1217 120 -1183
rect 60 -1251 120 -1217
rect 60 -1285 73 -1251
rect 107 -1285 120 -1251
rect 300 -1158 500 -1150
rect 300 -1170 349 -1158
rect 300 -1260 310 -1170
rect 383 -1192 417 -1158
rect 451 -1192 500 -1158
rect 350 -1210 500 -1192
rect 350 -1260 360 -1210
rect 300 -1270 360 -1260
rect 60 -1319 120 -1285
rect 60 -1353 73 -1319
rect 107 -1353 120 -1319
rect 60 -1387 120 -1353
rect 60 -1421 73 -1387
rect 107 -1421 120 -1387
rect 60 -1455 120 -1421
rect 60 -1489 73 -1455
rect 107 -1489 120 -1455
rect 60 -1523 120 -1489
rect 60 -1557 73 -1523
rect 107 -1557 120 -1523
rect 60 -1591 120 -1557
rect 800 -1500 870 -1067
rect 1000 -1123 1050 -1011
rect 1290 -909 1510 -860
rect 1290 -943 1293 -909
rect 1327 -943 1383 -909
rect 1417 -943 1471 -909
rect 1505 -943 1510 -909
rect 1290 -977 1510 -943
rect 1290 -1011 1293 -977
rect 1327 -1011 1383 -977
rect 1417 -1011 1471 -977
rect 1505 -1011 1510 -977
rect 1290 -1060 1510 -1011
rect 1740 -909 1790 -860
rect 1740 -943 1743 -909
rect 1777 -943 1790 -909
rect 1740 -977 1790 -943
rect 1740 -1011 1743 -977
rect 1777 -1011 1790 -977
rect 1000 -1157 1093 -1123
rect 1127 -1157 1143 -1123
rect 1740 -1130 1790 -1011
rect 1860 -909 1910 -810
rect 1860 -943 1873 -909
rect 1907 -943 1910 -909
rect 1860 -977 1910 -943
rect 1860 -1011 1873 -977
rect 1907 -1011 1910 -977
rect 1860 -1060 1910 -1011
rect 2030 -909 2090 -860
rect 2030 -943 2043 -909
rect 2077 -943 2090 -909
rect 2160 -910 2200 -810
rect 2030 -977 2090 -943
rect 2030 -1011 2043 -977
rect 2077 -1011 2090 -977
rect 2030 -1060 2090 -1011
rect 1912 -1130 1928 -1123
rect 1633 -1153 1667 -1137
rect 1000 -1299 1050 -1157
rect 1740 -1157 1928 -1130
rect 1962 -1130 1978 -1123
rect 1962 -1157 1980 -1130
rect 1740 -1170 1980 -1157
rect 1000 -1333 1013 -1299
rect 1047 -1333 1050 -1299
rect 1000 -1367 1050 -1333
rect 1000 -1401 1013 -1367
rect 1047 -1401 1050 -1367
rect 1000 -1450 1050 -1401
rect 1120 -1299 1170 -1250
rect 1120 -1333 1123 -1299
rect 1157 -1333 1170 -1299
rect 1120 -1340 1170 -1333
rect 1620 -1299 1670 -1250
rect 1620 -1333 1633 -1299
rect 1667 -1333 1670 -1299
rect 1620 -1340 1670 -1333
rect 1120 -1358 1670 -1340
rect 1120 -1367 1358 -1358
rect 1120 -1401 1123 -1367
rect 1157 -1392 1358 -1367
rect 1392 -1367 1670 -1358
rect 1392 -1392 1633 -1367
rect 1157 -1400 1633 -1392
rect 1157 -1401 1170 -1400
rect 1120 -1450 1170 -1401
rect 1620 -1401 1633 -1400
rect 1667 -1401 1670 -1367
rect 1240 -1468 1310 -1440
rect 1620 -1450 1670 -1401
rect 1740 -1299 1790 -1170
rect 2040 -1193 2090 -1060
rect 2150 -959 2200 -910
rect 2150 -993 2166 -959
rect 2150 -1027 2200 -993
rect 2150 -1061 2166 -1027
rect 2150 -1110 2200 -1061
rect 2280 -959 2340 -910
rect 2280 -993 2283 -959
rect 2317 -993 2340 -959
rect 2280 -1027 2340 -993
rect 2280 -1061 2283 -1027
rect 2317 -1061 2340 -1027
rect 2040 -1227 2043 -1193
rect 2077 -1227 2090 -1193
rect 2040 -1290 2090 -1227
rect 2280 -1203 2340 -1061
rect 2280 -1237 2293 -1203
rect 2327 -1237 2340 -1203
rect 1740 -1333 1743 -1299
rect 1777 -1333 1790 -1299
rect 1740 -1367 1790 -1333
rect 1740 -1401 1743 -1367
rect 1777 -1401 1790 -1367
rect 1870 -1320 2090 -1290
rect 2150 -1299 2210 -1250
rect 1870 -1343 2070 -1320
rect 1870 -1377 1919 -1343
rect 1953 -1377 1987 -1343
rect 2021 -1377 2070 -1343
rect 1870 -1380 2070 -1377
rect 2150 -1333 2173 -1299
rect 2207 -1333 2210 -1299
rect 2150 -1367 2210 -1333
rect 1740 -1450 1790 -1401
rect 2150 -1401 2173 -1367
rect 2207 -1401 2210 -1367
rect 800 -1513 1120 -1500
rect 800 -1547 1068 -1513
rect 1102 -1547 1120 -1513
rect 800 -1570 1120 -1547
rect 1240 -1523 1253 -1468
rect 1287 -1523 1310 -1468
rect 1780 -1520 1840 -1510
rect 1240 -1557 1310 -1523
rect 60 -1625 73 -1591
rect 107 -1625 120 -1591
rect 1240 -1591 1253 -1557
rect 1287 -1591 1310 -1557
rect 1240 -1620 1310 -1591
rect 1770 -1538 1840 -1520
rect 1770 -1572 1788 -1538
rect 1822 -1548 1840 -1538
rect 1770 -1582 1793 -1572
rect 1827 -1582 1840 -1548
rect 1770 -1610 1840 -1582
rect 60 -1659 120 -1625
rect 1880 -1623 2070 -1610
rect 60 -1693 73 -1659
rect 107 -1693 120 -1659
rect 1350 -1643 1500 -1640
rect 1350 -1677 1372 -1643
rect 1407 -1677 1444 -1643
rect 1478 -1677 1500 -1643
rect 1350 -1690 1500 -1677
rect 1880 -1657 1924 -1623
rect 1958 -1643 1992 -1623
rect 2026 -1640 2070 -1623
rect 2026 -1643 2080 -1640
rect 1961 -1657 1992 -1643
rect 1880 -1677 1927 -1657
rect 1961 -1677 1999 -1657
rect 2033 -1677 2080 -1643
rect 1880 -1690 2080 -1677
rect 2150 -1643 2210 -1401
rect 2280 -1299 2340 -1237
rect 2280 -1333 2288 -1299
rect 2322 -1333 2340 -1299
rect 2280 -1367 2340 -1333
rect 2280 -1401 2288 -1367
rect 2322 -1401 2340 -1367
rect 2280 -1450 2340 -1401
rect 2150 -1677 2163 -1643
rect 2197 -1677 2210 -1643
rect 2150 -1690 2210 -1677
rect 60 -1727 120 -1693
rect 60 -1761 73 -1727
rect 107 -1761 120 -1727
rect 60 -1795 120 -1761
rect 60 -1829 73 -1795
rect 107 -1829 120 -1795
rect 60 -1863 120 -1829
rect 60 -1897 73 -1863
rect 107 -1897 120 -1863
rect 60 -1931 120 -1897
rect 60 -1965 73 -1931
rect 107 -1965 120 -1931
rect 60 -1999 120 -1965
rect 60 -2033 73 -1999
rect 107 -2033 120 -1999
rect 60 -2067 120 -2033
rect 60 -2101 73 -2067
rect 107 -2101 120 -2067
rect 60 -2135 120 -2101
rect 60 -2169 73 -2135
rect 107 -2169 120 -2135
rect -150 -2188 -60 -2180
rect -150 -2222 -122 -2188
rect -88 -2222 -60 -2188
rect -150 -2268 -60 -2222
rect -150 -2302 -122 -2268
rect -88 -2302 -60 -2268
rect -150 -2330 -60 -2302
rect 60 -2250 120 -2169
rect 250 -2170 310 -2164
rect 240 -2193 470 -2170
rect 240 -2227 263 -2193
rect 297 -2227 413 -2193
rect 447 -2227 470 -2193
rect 240 -2250 470 -2227
rect 60 -2320 110 -2250
rect 250 -2256 310 -2250
rect -20 -2360 110 -2320
rect -20 -2400 30 -2360
rect 447 -2382 463 -2348
rect 497 -2382 513 -2348
rect -30 -2430 30 -2400
rect -30 -2464 -17 -2430
rect 17 -2464 30 -2430
rect -30 -2498 30 -2464
rect -30 -2532 -17 -2498
rect 17 -2532 30 -2498
rect -30 -2566 30 -2532
rect -30 -2600 -17 -2566
rect 17 -2600 30 -2566
rect -30 -2640 30 -2600
rect 250 -2430 390 -2400
rect 250 -2464 263 -2430
rect 297 -2435 390 -2430
rect 297 -2464 343 -2435
rect 250 -2469 343 -2464
rect 377 -2469 390 -2435
rect 250 -2498 390 -2469
rect 250 -2532 263 -2498
rect 297 -2503 390 -2498
rect 297 -2532 343 -2503
rect 250 -2537 343 -2532
rect 377 -2537 390 -2503
rect 250 -2540 390 -2537
rect 250 -2566 520 -2540
rect 250 -2600 263 -2566
rect 297 -2571 520 -2566
rect 297 -2600 343 -2571
rect 250 -2605 343 -2600
rect 377 -2573 520 -2571
rect 377 -2605 402 -2573
rect 250 -2607 402 -2605
rect 436 -2607 474 -2573
rect 508 -2607 520 -2573
rect 250 -2640 520 -2607
<< viali >>
rect 923 218 957 252
rect 2653 223 2687 257
rect 1183 -197 1217 -163
rect 2473 -107 2497 -78
rect 2497 -107 2507 -78
rect 2473 -112 2507 -107
rect 2038 -197 2072 -163
rect 8 -417 42 -383
rect 537 -427 571 -393
rect 609 -427 643 -393
rect 517 -767 539 -743
rect 539 -767 551 -743
rect 589 -767 607 -743
rect 607 -767 623 -743
rect 2658 -398 2692 -388
rect 2658 -422 2692 -398
rect 2643 -667 2677 -633
rect 517 -777 551 -767
rect 589 -777 623 -767
rect 1179 -792 1213 -758
rect 1251 -792 1285 -758
rect 1323 -792 1357 -758
rect 1395 -792 1429 -758
rect 1467 -792 1501 -758
rect 1539 -792 1573 -758
rect 1611 -792 1645 -758
rect 1683 -792 1717 -758
rect 1755 -792 1789 -758
rect 1827 -792 1861 -758
rect 1899 -792 1933 -758
rect 1971 -792 2005 -758
rect 2043 -792 2077 -758
rect 2115 -792 2149 -758
rect 2187 -792 2221 -758
rect -147 -937 -113 -903
rect 593 -997 627 -963
rect 818 -1067 852 -1033
rect 310 -1192 349 -1170
rect 349 -1192 350 -1170
rect 310 -1260 350 -1192
rect 1633 -1187 1667 -1178
rect 1633 -1212 1667 -1187
rect 2293 -1237 2327 -1203
rect 1068 -1547 1102 -1513
rect 1253 -1489 1287 -1468
rect 1253 -1502 1287 -1489
rect 1788 -1548 1822 -1538
rect 1788 -1572 1793 -1548
rect 1793 -1572 1822 -1548
rect 1372 -1677 1373 -1643
rect 1373 -1677 1406 -1643
rect 1444 -1677 1478 -1643
rect 1927 -1657 1958 -1643
rect 1958 -1657 1961 -1643
rect 1999 -1657 2026 -1643
rect 2026 -1657 2033 -1643
rect 1927 -1677 1961 -1657
rect 1999 -1677 2033 -1657
rect 2163 -1677 2197 -1643
rect -122 -2222 -88 -2188
rect 413 -2227 447 -2193
rect 463 -2382 497 -2348
rect 402 -2607 436 -2573
rect 474 -2607 508 -2573
<< metal1 >>
rect -200 257 2800 270
rect -200 252 2653 257
rect -200 218 923 252
rect 957 223 2653 252
rect 2687 223 2800 257
rect 957 218 2800 223
rect -200 120 2800 218
rect -16 -365 66 -353
rect -16 -383 185 -365
rect -16 -417 8 -383
rect 42 -417 185 -383
rect -16 -435 185 -417
rect -16 -447 66 -435
rect 115 -615 185 -435
rect 490 -380 590 120
rect 2440 -74 2540 -50
rect 2440 -78 2534 -74
rect 2440 -112 2473 -78
rect 2507 -112 2534 -78
rect 2440 -126 2534 -112
rect 2586 -126 2592 -74
rect 2440 -140 2540 -126
rect 1174 -150 1226 -148
rect 644 -154 1230 -150
rect 644 -206 654 -154
rect 706 -163 1232 -154
rect 706 -197 1183 -163
rect 1217 -197 1232 -163
rect 706 -206 1232 -197
rect 2018 -163 2092 -149
rect 2018 -197 2038 -163
rect 2072 -197 2092 -163
rect 644 -210 1230 -206
rect 1174 -212 1226 -210
rect 2018 -211 2092 -197
rect 490 -393 690 -380
rect 490 -427 537 -393
rect 571 -427 609 -393
rect 643 -427 690 -393
rect 2030 -423 2080 -211
rect 490 -440 690 -427
rect 735 -473 2080 -423
rect 2640 -388 2710 -360
rect 2640 -422 2658 -388
rect 2692 -422 2710 -388
rect 2640 -449 2710 -422
rect 109 -624 191 -615
rect 109 -676 124 -624
rect 176 -676 191 -624
rect 109 -685 191 -676
rect 115 -730 185 -685
rect 510 -730 650 -720
rect 490 -734 650 -730
rect 490 -786 512 -734
rect 564 -786 576 -734
rect 628 -786 650 -734
rect 490 -790 650 -786
rect 490 -810 640 -790
rect 735 -855 785 -473
rect 2640 -501 2649 -449
rect 2701 -501 2710 -449
rect 2640 -516 2710 -501
rect 2630 -620 2690 -614
rect 2624 -624 2696 -620
rect 2624 -676 2634 -624
rect 2686 -676 2696 -624
rect 2624 -680 2696 -676
rect 2630 -686 2690 -680
rect 970 -758 2290 -730
rect 860 -770 920 -764
rect 970 -770 1179 -758
rect 860 -774 1179 -770
rect 860 -826 864 -774
rect 916 -792 1179 -774
rect 1213 -792 1251 -758
rect 1285 -792 1323 -758
rect 1357 -792 1395 -758
rect 1429 -792 1467 -758
rect 1501 -792 1539 -758
rect 1573 -792 1611 -758
rect 1645 -792 1683 -758
rect 1717 -792 1755 -758
rect 1789 -792 1827 -758
rect 1861 -792 1899 -758
rect 1933 -792 1971 -758
rect 2005 -792 2043 -758
rect 2077 -792 2115 -758
rect 2149 -792 2187 -758
rect 2221 -770 2290 -758
rect 2221 -774 2626 -770
rect 2221 -792 2564 -774
rect 916 -826 2564 -792
rect 2616 -826 2626 -774
rect 860 -830 2626 -826
rect 860 -836 920 -830
rect -153 -903 -107 -891
rect -22 -903 -16 -894
rect -153 -937 -147 -903
rect -113 -937 -16 -903
rect -153 -949 -107 -937
rect -22 -946 -16 -937
rect 36 -946 42 -894
rect 300 -905 785 -855
rect 300 -1150 340 -905
rect 584 -954 636 -948
rect 578 -1006 584 -954
rect 636 -1006 642 -954
rect 584 -1012 636 -1006
rect 794 -1009 876 -1003
rect 788 -1024 876 -1009
rect 788 -1076 803 -1024
rect 855 -1076 876 -1024
rect 788 -1091 876 -1076
rect 794 -1097 876 -1091
rect 300 -1170 360 -1150
rect 300 -1260 310 -1170
rect 350 -1260 360 -1170
rect 1624 -1169 1676 -1163
rect 2274 -1180 2346 -1178
rect 1624 -1227 1676 -1221
rect 2270 -1199 2390 -1180
rect 2270 -1203 2314 -1199
rect 2270 -1237 2293 -1203
rect 414 -1254 466 -1248
rect 300 -1300 414 -1260
rect 2270 -1251 2314 -1237
rect 2366 -1251 2390 -1199
rect 2270 -1270 2390 -1251
rect 414 -1312 466 -1306
rect -470 -1410 3090 -1350
rect 1230 -1468 1310 -1440
rect 1230 -1488 1253 -1468
rect 1214 -1494 1253 -1488
rect 1062 -1504 1108 -1501
rect 1287 -1502 1310 -1468
rect 1053 -1556 1059 -1504
rect 1111 -1556 1117 -1504
rect 1266 -1530 1310 -1502
rect 1760 -1510 1790 -1410
rect 1760 -1520 1840 -1510
rect 1214 -1552 1266 -1546
rect 1760 -1538 1850 -1520
rect 1062 -1559 1108 -1556
rect 1760 -1572 1788 -1538
rect 1822 -1572 1850 -1538
rect 1760 -1590 1850 -1572
rect 635 -1625 705 -1615
rect 635 -1643 2330 -1625
rect 635 -1677 1372 -1643
rect 1406 -1677 1444 -1643
rect 1478 -1677 1927 -1643
rect 1961 -1677 1999 -1643
rect 2033 -1677 2163 -1643
rect 2197 -1677 2330 -1643
rect 635 -1695 2330 -1677
rect -150 -2109 -60 -2090
rect -150 -2161 -131 -2109
rect -79 -2161 -60 -2109
rect -150 -2188 -60 -2161
rect 384 -2164 476 -2158
rect -150 -2222 -122 -2188
rect -88 -2222 -60 -2188
rect -150 -2240 -60 -2222
rect 378 -2178 482 -2164
rect 378 -2230 404 -2178
rect 456 -2230 482 -2178
rect 378 -2256 482 -2230
rect 454 -2339 506 -2333
rect 451 -2388 454 -2342
rect 506 -2388 509 -2342
rect 454 -2397 506 -2391
rect 635 -2520 705 -1695
rect -200 -2544 2800 -2520
rect -200 -2573 564 -2544
rect -200 -2607 402 -2573
rect 436 -2607 474 -2573
rect 508 -2596 564 -2573
rect 616 -2594 2800 -2544
rect 616 -2596 2569 -2594
rect 508 -2607 2569 -2596
rect -200 -2646 2569 -2607
rect 2621 -2646 2800 -2594
rect -200 -2670 2800 -2646
<< via1 >>
rect 2534 -126 2586 -74
rect 654 -206 706 -154
rect 124 -676 176 -624
rect 512 -743 564 -734
rect 512 -777 517 -743
rect 517 -777 551 -743
rect 551 -777 564 -743
rect 512 -786 564 -777
rect 576 -743 628 -734
rect 576 -777 589 -743
rect 589 -777 623 -743
rect 623 -777 628 -743
rect 576 -786 628 -777
rect 2649 -501 2701 -449
rect 2634 -633 2686 -624
rect 2634 -667 2643 -633
rect 2643 -667 2677 -633
rect 2677 -667 2686 -633
rect 2634 -676 2686 -667
rect 864 -826 916 -774
rect 2564 -826 2616 -774
rect -16 -946 36 -894
rect 584 -963 636 -954
rect 584 -997 593 -963
rect 593 -997 627 -963
rect 627 -997 636 -963
rect 584 -1006 636 -997
rect 803 -1033 855 -1024
rect 803 -1067 818 -1033
rect 818 -1067 852 -1033
rect 852 -1067 855 -1033
rect 803 -1076 855 -1067
rect 1624 -1178 1676 -1169
rect 1624 -1212 1633 -1178
rect 1633 -1212 1667 -1178
rect 1667 -1212 1676 -1178
rect 1624 -1221 1676 -1212
rect 2314 -1203 2366 -1199
rect 2314 -1237 2327 -1203
rect 2327 -1237 2366 -1203
rect 414 -1306 466 -1254
rect 2314 -1251 2366 -1237
rect 1214 -1502 1253 -1494
rect 1253 -1502 1266 -1494
rect 1059 -1513 1111 -1504
rect 1059 -1547 1068 -1513
rect 1068 -1547 1102 -1513
rect 1102 -1547 1111 -1513
rect 1059 -1556 1111 -1547
rect 1214 -1546 1266 -1502
rect -131 -2161 -79 -2109
rect 404 -2193 456 -2178
rect 404 -2227 413 -2193
rect 413 -2227 447 -2193
rect 447 -2227 456 -2193
rect 404 -2230 456 -2227
rect 454 -2348 506 -2339
rect 454 -2382 463 -2348
rect 463 -2382 497 -2348
rect 497 -2382 506 -2348
rect 454 -2391 506 -2382
rect 564 -2596 616 -2544
rect 2569 -2646 2621 -2594
<< metal2 >>
rect -140 -2109 -70 570
rect -10 -888 60 570
rect 115 -610 185 -609
rect 110 -622 190 -610
rect 110 -678 122 -622
rect 178 -678 190 -622
rect 110 -690 190 -678
rect 115 -691 185 -690
rect -16 -894 60 -888
rect 36 -903 60 -894
rect 36 -937 77 -903
rect 36 -946 60 -937
rect -16 -952 60 -946
rect -140 -2161 -131 -2109
rect -79 -2161 -70 -2109
rect -140 -2730 -70 -2161
rect -10 -2950 60 -952
rect 220 -960 290 570
rect 650 -150 710 -144
rect 641 -152 719 -150
rect 641 -208 652 -152
rect 708 -208 719 -152
rect 641 -210 719 -208
rect 650 -216 710 -210
rect 939 -685 969 570
rect 1104 -640 1144 570
rect 939 -715 1005 -685
rect 1104 -690 1180 -640
rect 475 -723 780 -715
rect 475 -734 805 -723
rect 475 -786 512 -734
rect 564 -786 576 -734
rect 628 -786 805 -734
rect 475 -825 805 -786
rect 670 -865 805 -825
rect 850 -772 930 -760
rect 850 -828 862 -772
rect 918 -828 930 -772
rect 850 -840 930 -828
rect 584 -954 636 -948
rect 220 -1000 584 -960
rect 220 -2785 290 -1000
rect 666 -965 805 -865
rect 975 -885 1005 -715
rect 584 -1012 636 -1006
rect 670 -990 805 -965
rect 939 -915 1005 -885
rect 670 -1024 870 -990
rect 670 -1076 803 -1024
rect 855 -1076 870 -1024
rect 670 -1210 870 -1076
rect 670 -1215 805 -1210
rect 408 -1306 414 -1254
rect 466 -1260 472 -1254
rect 466 -1300 610 -1260
rect 466 -1306 472 -1300
rect 384 -2164 476 -2155
rect 378 -2176 482 -2164
rect 378 -2232 402 -2176
rect 458 -2232 482 -2176
rect 378 -2244 482 -2232
rect 384 -2253 476 -2244
rect 450 -2337 510 -2326
rect 450 -2339 452 -2337
rect 508 -2339 510 -2337
rect 448 -2391 452 -2339
rect 508 -2391 512 -2339
rect 450 -2393 452 -2391
rect 508 -2393 510 -2391
rect 450 -2404 510 -2393
rect 570 -2544 610 -1300
rect 670 -1318 794 -1215
rect 661 -1352 803 -1318
rect 661 -1408 704 -1352
rect 760 -1408 803 -1352
rect 661 -1442 803 -1408
rect 939 -1735 969 -915
rect 1059 -1504 1111 -1498
rect 1059 -1562 1111 -1556
rect 1140 -1630 1180 -690
rect 1210 -1492 1270 -1481
rect 1210 -1494 1212 -1492
rect 1268 -1494 1270 -1492
rect 1208 -1546 1212 -1494
rect 1268 -1546 1272 -1494
rect 1210 -1548 1212 -1546
rect 1268 -1548 1270 -1546
rect 1210 -1559 1270 -1548
rect 1104 -1670 1180 -1630
rect 1104 -1730 1144 -1670
rect 1374 -1735 1404 570
rect 1539 -1730 1579 570
rect 1610 -922 1690 -901
rect 1610 -978 1622 -922
rect 1678 -978 1690 -922
rect 1610 -1169 1690 -978
rect 1610 -1221 1624 -1169
rect 1676 -1221 1690 -1169
rect 1610 -1240 1690 -1221
rect 1809 -1725 1839 570
rect 1974 -1740 2014 570
rect 2244 -805 2274 570
rect 2236 -806 2274 -805
rect 2205 -835 2274 -806
rect 2205 -1345 2235 -835
rect 2409 -1040 2449 570
rect 2530 48 2590 59
rect 2530 -8 2532 48
rect 2588 -8 2590 48
rect 2530 -19 2590 -8
rect 2540 -68 2580 -19
rect 2534 -74 2586 -68
rect 2534 -132 2586 -126
rect 2640 -440 2710 -431
rect 2634 -447 2716 -440
rect 2634 -503 2647 -447
rect 2703 -503 2716 -447
rect 2634 -510 2716 -503
rect 2640 -519 2710 -510
rect 2632 -620 2688 -613
rect 2624 -622 2696 -620
rect 2624 -678 2632 -622
rect 2688 -678 2696 -622
rect 2624 -680 2696 -678
rect 2632 -687 2688 -680
rect 2560 -770 2620 -764
rect 2551 -772 2629 -770
rect 2551 -828 2562 -772
rect 2618 -828 2629 -772
rect 2551 -830 2629 -828
rect 2560 -836 2620 -830
rect 2410 -1060 2449 -1040
rect 2410 -1100 2510 -1060
rect 2300 -1197 2390 -1180
rect 2300 -1253 2312 -1197
rect 2368 -1253 2390 -1197
rect 2300 -1270 2390 -1253
rect 2470 -1310 2510 -1100
rect 2205 -1375 2274 -1345
rect 2244 -1735 2274 -1375
rect 2409 -1350 2510 -1310
rect 2409 -1700 2449 -1350
rect 558 -2596 564 -2544
rect 616 -2596 622 -2544
rect 939 -2935 969 -2450
rect 1104 -2940 1144 -2430
rect 1374 -2940 1404 -2445
rect 1539 -2940 1579 -2440
rect 1809 -2940 1839 -2445
rect 1974 -2940 2014 -2440
rect 2244 -2940 2274 -2445
rect 2409 -2940 2449 -2440
rect 2560 -2585 2630 -1730
rect 2554 -2594 2636 -2585
rect 2554 -2646 2569 -2594
rect 2621 -2646 2636 -2594
rect 2554 -2655 2636 -2646
<< via2 >>
rect 122 -624 178 -622
rect 122 -676 124 -624
rect 124 -676 176 -624
rect 176 -676 178 -624
rect 122 -678 178 -676
rect 652 -154 708 -152
rect 652 -206 654 -154
rect 654 -206 706 -154
rect 706 -206 708 -154
rect 652 -208 708 -206
rect 862 -774 918 -772
rect 862 -826 864 -774
rect 864 -826 916 -774
rect 916 -826 918 -774
rect 862 -828 918 -826
rect 402 -2178 458 -2176
rect 402 -2230 404 -2178
rect 404 -2230 456 -2178
rect 456 -2230 458 -2178
rect 402 -2232 458 -2230
rect 452 -2339 508 -2337
rect 452 -2391 454 -2339
rect 454 -2391 506 -2339
rect 506 -2391 508 -2339
rect 452 -2393 508 -2391
rect 704 -1408 760 -1352
rect 1212 -1494 1268 -1492
rect 1212 -1546 1214 -1494
rect 1214 -1546 1266 -1494
rect 1266 -1546 1268 -1494
rect 1212 -1548 1268 -1546
rect 1622 -978 1678 -922
rect 2532 -8 2588 48
rect 2647 -449 2703 -447
rect 2647 -501 2649 -449
rect 2649 -501 2701 -449
rect 2701 -501 2703 -449
rect 2647 -503 2703 -501
rect 2632 -624 2688 -622
rect 2632 -676 2634 -624
rect 2634 -676 2686 -624
rect 2686 -676 2688 -624
rect 2632 -678 2688 -676
rect 2562 -774 2618 -772
rect 2562 -826 2564 -774
rect 2564 -826 2616 -774
rect 2616 -826 2618 -774
rect 2562 -828 2618 -826
rect 2312 -1199 2368 -1197
rect 2312 -1251 2314 -1199
rect 2314 -1251 2366 -1199
rect 2366 -1251 2368 -1199
rect 2312 -1253 2368 -1251
<< metal3 >>
rect 2525 50 2595 55
rect -300 48 3090 50
rect -300 -8 2532 48
rect 2588 -8 3090 48
rect -300 -10 3090 -8
rect 2525 -15 2595 -10
rect 645 -150 715 -145
rect -470 -152 3090 -150
rect -470 -208 652 -152
rect 708 -208 3090 -152
rect -470 -210 3090 -208
rect 645 -215 715 -210
rect 2635 -447 2715 -435
rect 2635 -450 2647 -447
rect -370 -503 2647 -450
rect 2703 -450 2715 -447
rect 2703 -503 3050 -450
rect -370 -510 3050 -503
rect 2635 -515 2715 -510
rect 100 -618 200 -600
rect 2640 -617 2780 -590
rect 100 -682 118 -618
rect 182 -682 200 -618
rect 100 -700 200 -682
rect 2627 -618 2780 -617
rect 2627 -622 2701 -618
rect 2627 -678 2632 -622
rect 2688 -678 2701 -622
rect 2627 -682 2701 -678
rect 2765 -682 2780 -618
rect 2627 -683 2780 -682
rect 2640 -700 2780 -683
rect 857 -770 923 -767
rect 2555 -770 2625 -765
rect -450 -772 923 -770
rect -450 -828 862 -772
rect 918 -828 923 -772
rect -450 -830 923 -828
rect 2350 -772 3090 -770
rect 2350 -828 2562 -772
rect 2618 -828 3090 -772
rect 2350 -830 3090 -828
rect 857 -833 923 -830
rect 2555 -835 2625 -830
rect -370 -922 3090 -900
rect -370 -960 1622 -922
rect 1605 -978 1622 -960
rect 1678 -960 3090 -922
rect 1678 -978 1695 -960
rect 1605 -995 1695 -978
rect -340 -1130 3090 -1070
rect 100 -1318 560 -1310
rect 665 -1318 799 -1313
rect 100 -1352 799 -1318
rect 100 -1408 704 -1352
rect 760 -1408 799 -1352
rect 100 -1442 799 -1408
rect 100 -1770 560 -1442
rect 665 -1447 799 -1442
rect 1210 -1485 1270 -1130
rect 2305 -1197 2539 -1190
rect 2305 -1253 2312 -1197
rect 2368 -1253 2539 -1197
rect 2305 -1260 2539 -1253
rect 1205 -1492 1275 -1485
rect 1205 -1548 1212 -1492
rect 1268 -1548 1275 -1492
rect 1205 -1555 1275 -1548
rect 2479 -1790 2539 -1260
rect 130 -2040 680 -2030
rect 120 -2090 680 -2040
rect 120 -2260 180 -2090
rect 379 -2167 481 -2153
rect 379 -2231 398 -2167
rect 462 -2231 481 -2167
rect 379 -2232 402 -2231
rect 458 -2232 481 -2231
rect 379 -2249 481 -2232
rect -470 -2320 180 -2260
rect 620 -2260 680 -2090
rect 620 -2320 3080 -2260
rect 430 -2337 520 -2330
rect 430 -2393 452 -2337
rect 508 -2393 520 -2337
rect 430 -2520 520 -2393
rect -200 -2580 3090 -2520
<< via3 >>
rect 118 -622 182 -618
rect 118 -678 122 -622
rect 122 -678 178 -622
rect 178 -678 182 -622
rect 118 -682 182 -678
rect 2701 -682 2765 -618
rect 398 -2176 462 -2167
rect 398 -2231 402 -2176
rect 402 -2231 458 -2176
rect 458 -2231 462 -2176
<< mimcap >>
rect 130 -1422 530 -1340
rect 130 -1646 361 -1422
rect 505 -1646 530 -1422
rect 130 -1740 530 -1646
<< mimcapcontact >>
rect 361 -1646 505 -1422
<< metal4 >>
rect 115 -618 185 -615
rect 115 -682 118 -618
rect 182 -682 185 -618
rect 115 -1029 185 -682
rect 109 -1101 191 -1029
rect 115 -1195 185 -1101
rect 270 -1195 670 -1190
rect 115 -1239 670 -1195
rect 115 -1265 704 -1239
rect 270 -1422 704 -1265
rect 270 -1646 361 -1422
rect 505 -1646 704 -1422
rect 270 -1740 704 -1646
rect 349 -1802 704 -1740
rect 349 -1849 412 -1802
rect 350 -1850 412 -1849
rect 370 -2038 412 -1850
rect 648 -1849 704 -1802
rect 648 -2038 690 -1849
rect 370 -2080 690 -2038
rect 390 -2158 470 -2080
rect 378 -2167 482 -2158
rect 378 -2231 398 -2167
rect 462 -2231 482 -2167
rect 378 -2240 482 -2231
rect 814 -2940 874 570
rect 1004 -1740 1064 570
rect 1249 -1740 1309 570
rect 1439 -1740 1499 570
rect 1684 -1740 1744 570
rect 1874 -1740 1934 570
rect 2119 -1740 2179 570
rect 2309 -1740 2369 570
rect 2700 -618 2800 570
rect 2700 -682 2701 -618
rect 2765 -682 2800 -618
rect 1004 -2930 1064 -2400
rect 1249 -2940 1309 -2420
rect 1439 -2940 1499 -2420
rect 1684 -2940 1744 -2420
rect 1874 -2940 1934 -2420
rect 2119 -2940 2179 -2420
rect 2309 -2940 2369 -2420
rect 2560 -2645 2630 -1730
rect 2700 -3000 2800 -682
<< via4 >>
rect 412 -2038 648 -1802
<< metal5 >>
rect -360 140 2960 460
rect -360 -2540 -40 140
rect 280 -1802 2320 -180
rect 280 -2038 412 -1802
rect 648 -2038 2320 -1802
rect 280 -2220 2320 -2038
rect 2640 -2540 2960 140
rect -360 -2860 2960 -2540
<< glass >>
rect 480 -2020 2120 -380
use 8bit_dram  8bit_dram_0 ~/topmetal_dps/magic/ram
timestamp 1661550438
transform -1 0 2469 0 -1 -1700
box -70 -20 1745 780
<< labels >>
rlabel poly s 2150 -70 2150 -70 4 AMP_OUT
port 1 nsew
rlabel metal5 s 2700 -1680 2700 -1680 4 gring
port 2 nsew
rlabel metal1 s -170 240 -170 240 4 VDD
port 3 nsew
rlabel metal2 s -130 260 -130 260 4 VREF
port 4 nsew
rlabel metal4 s 2730 510 2730 510 4 PIX_OUT
port 5 nsew
rlabel metal3 s 3020 -480 3020 -480 4 ROW_SEL
port 6 nsew
rlabel metal3 s 3020 -180 3020 -180 4 CSA_VREF
port 7 nsew
rlabel metal3 s 3040 20 3040 20 4 SF_IB
port 8 nsew
rlabel metal3 s 3060 -2560 3060 -2560 4 NB1
port 9 nsew
rlabel metal1 s 2630 -2620 2630 -2620 4 GND
port 10 nsew
rlabel metal3 s 3020 -800 3020 -800 4 DVDD
port 11 nsew
rlabel metal5 s 352 -1964 352 -1964 4 PIX_IN
port 12 nsew
rlabel metal3 s 3022 -2286 3022 -2286 4 READ
port 13 nsew
rlabel metal1 s 3022 -1382 3022 -1382 4 BIAS2
port 14 nsew
rlabel metal3 s 3027 -1112 3027 -1112 4 BIAS1
port 15 nsew
rlabel metal3 s 2999 -929 2999 -929 4 V_RAMP
port 16 nsew
rlabel metal2 s 2431 -2902 2431 -2902 4 GRAYx0x
port 17 nsew
rlabel metal2 s 2256 -2915 2256 -2915 4 OUTx1x
port 18 nsew
rlabel metal4 s 2135 -2917 2135 -2917 4 OUTx0x
port 19 nsew
rlabel metal2 s 1821 -2906 1821 -2906 4 OUTx3x
port 20 nsew
rlabel metal4 s 1716 -2898 1716 -2898 4 OUTx2x
port 21 nsew
rlabel metal2 s 1388 -2908 1388 -2908 4 OUTx5x
port 22 nsew
rlabel metal4 s 1283 -2898 1283 -2898 4 OUTx4x
port 23 nsew
rlabel metal2 s 1119 -2906 1119 -2906 4 GRAYx6x
port 24 nsew
rlabel metal4 s 1031 -2900 1031 -2900 4 GRAYx7x
port 25 nsew
rlabel metal4 s 841 -2921 841 -2921 4 OUTx6x
port 26 nsew
rlabel metal2 s 959 -2895 959 -2895 4 OUTx7x
port 27 nsew
rlabel metal4 s 1470 -2910 1470 -2910 4 GRAYx5x
port 28 nsew
rlabel metal2 s 1553 -2891 1553 -2891 4 GRAYx4x
port 29 nsew
rlabel metal4 s 1903 -2922 1903 -2922 4 GRAYx3x
port 30 nsew
rlabel metal2 s 1989 -2907 1989 -2907 4 GRAYx2x
port 31 nsew
rlabel metal4 s 2341 -2908 2341 -2908 4 GRAYx1x
port 32 nsew
rlabel metal2 s 20 510 20 510 4 VBIAS
port 33 nsew
rlabel metal2 s 270 520 270 520 4 NB2
port 34 nsew
<< end >>
