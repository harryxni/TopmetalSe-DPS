magic
tech sky130B
magscale 1 2
timestamp 1606063140
<< nwell >>
rect -992 -497 992 497
<< mvpmos >>
rect -734 -200 -574 200
rect -516 -200 -356 200
rect -298 -200 -138 200
rect -80 -200 80 200
rect 138 -200 298 200
rect 356 -200 516 200
rect 574 -200 734 200
<< mvpdiff >>
rect -792 188 -734 200
rect -792 -188 -780 188
rect -746 -188 -734 188
rect -792 -200 -734 -188
rect -574 188 -516 200
rect -574 -188 -562 188
rect -528 -188 -516 188
rect -574 -200 -516 -188
rect -356 188 -298 200
rect -356 -188 -344 188
rect -310 -188 -298 188
rect -356 -200 -298 -188
rect -138 188 -80 200
rect -138 -188 -126 188
rect -92 -188 -80 188
rect -138 -200 -80 -188
rect 80 188 138 200
rect 80 -188 92 188
rect 126 -188 138 188
rect 80 -200 138 -188
rect 298 188 356 200
rect 298 -188 310 188
rect 344 -188 356 188
rect 298 -200 356 -188
rect 516 188 574 200
rect 516 -188 528 188
rect 562 -188 574 188
rect 516 -200 574 -188
rect 734 188 792 200
rect 734 -188 746 188
rect 780 -188 792 188
rect 734 -200 792 -188
<< mvpdiffc >>
rect -780 -188 -746 188
rect -562 -188 -528 188
rect -344 -188 -310 188
rect -126 -188 -92 188
rect 92 -188 126 188
rect 310 -188 344 188
rect 528 -188 562 188
rect 746 -188 780 188
<< mvnsubdiff >>
rect -926 419 926 431
rect -926 385 -818 419
rect 818 385 926 419
rect -926 373 926 385
rect -926 323 -868 373
rect -926 -323 -914 323
rect -880 -323 -868 323
rect 868 323 926 373
rect -926 -373 -868 -323
rect 868 -323 880 323
rect 914 -323 926 323
rect 868 -373 926 -323
rect -926 -385 926 -373
rect -926 -419 -818 -385
rect 818 -419 926 -385
rect -926 -431 926 -419
<< mvnsubdiffcont >>
rect -818 385 818 419
rect -914 -323 -880 323
rect 880 -323 914 323
rect -818 -419 818 -385
<< poly >>
rect -734 281 -574 297
rect -734 247 -718 281
rect -590 247 -574 281
rect -734 200 -574 247
rect -516 281 -356 297
rect -516 247 -500 281
rect -372 247 -356 281
rect -516 200 -356 247
rect -298 281 -138 297
rect -298 247 -282 281
rect -154 247 -138 281
rect -298 200 -138 247
rect -80 281 80 297
rect -80 247 -64 281
rect 64 247 80 281
rect -80 200 80 247
rect 138 281 298 297
rect 138 247 154 281
rect 282 247 298 281
rect 138 200 298 247
rect 356 281 516 297
rect 356 247 372 281
rect 500 247 516 281
rect 356 200 516 247
rect 574 281 734 297
rect 574 247 590 281
rect 718 247 734 281
rect 574 200 734 247
rect -734 -247 -574 -200
rect -734 -281 -718 -247
rect -590 -281 -574 -247
rect -734 -297 -574 -281
rect -516 -247 -356 -200
rect -516 -281 -500 -247
rect -372 -281 -356 -247
rect -516 -297 -356 -281
rect -298 -247 -138 -200
rect -298 -281 -282 -247
rect -154 -281 -138 -247
rect -298 -297 -138 -281
rect -80 -247 80 -200
rect -80 -281 -64 -247
rect 64 -281 80 -247
rect -80 -297 80 -281
rect 138 -247 298 -200
rect 138 -281 154 -247
rect 282 -281 298 -247
rect 138 -297 298 -281
rect 356 -247 516 -200
rect 356 -281 372 -247
rect 500 -281 516 -247
rect 356 -297 516 -281
rect 574 -247 734 -200
rect 574 -281 590 -247
rect 718 -281 734 -247
rect 574 -297 734 -281
<< polycont >>
rect -718 247 -590 281
rect -500 247 -372 281
rect -282 247 -154 281
rect -64 247 64 281
rect 154 247 282 281
rect 372 247 500 281
rect 590 247 718 281
rect -718 -281 -590 -247
rect -500 -281 -372 -247
rect -282 -281 -154 -247
rect -64 -281 64 -247
rect 154 -281 282 -247
rect 372 -281 500 -247
rect 590 -281 718 -247
<< locali >>
rect -914 385 -818 419
rect 818 385 914 419
rect 880 323 914 385
rect -734 247 -718 281
rect -590 247 -574 281
rect -516 247 -500 281
rect -372 247 -356 281
rect -298 247 -282 281
rect -154 247 -138 281
rect -80 247 -64 281
rect 64 247 80 281
rect 138 247 154 281
rect 282 247 298 281
rect 356 247 372 281
rect 500 247 516 281
rect 574 247 590 281
rect 718 247 734 281
rect -780 188 -746 204
rect -780 -204 -746 -188
rect -562 188 -528 204
rect -562 -204 -528 -188
rect -344 188 -310 204
rect -344 -204 -310 -188
rect -126 188 -92 204
rect -126 -204 -92 -188
rect 92 188 126 204
rect 92 -204 126 -188
rect 310 188 344 204
rect 310 -204 344 -188
rect 528 188 562 204
rect 528 -204 562 -188
rect 746 188 780 204
rect 746 -204 780 -188
rect -734 -281 -718 -247
rect -590 -281 -574 -247
rect -516 -281 -500 -247
rect -372 -281 -356 -247
rect -298 -281 -282 -247
rect -154 -281 -138 -247
rect -80 -281 -64 -247
rect 64 -281 80 -247
rect 138 -281 154 -247
rect 282 -281 298 -247
rect 356 -281 372 -247
rect 500 -281 516 -247
rect 574 -281 590 -247
rect 718 -281 734 -247
rect -914 -385 -880 -323
rect 880 -385 914 -323
rect -914 -419 -818 -385
rect 818 -419 914 -385
<< viali >>
rect -792 385 792 419
rect -914 323 -880 385
rect -914 38 -880 323
rect -718 247 -590 281
rect -500 247 -372 281
rect -282 247 -154 281
rect -64 247 64 281
rect 154 247 282 281
rect 372 247 500 281
rect 590 247 718 281
rect -780 21 -746 171
rect -562 -171 -528 -21
rect -344 21 -310 171
rect -126 -171 -92 -21
rect 92 21 126 171
rect 310 -171 344 -21
rect 528 21 562 171
rect 746 -171 780 -21
rect -718 -281 -590 -247
rect -500 -281 -372 -247
rect -282 -281 -154 -247
rect -64 -281 64 -247
rect 154 -281 282 -247
rect 372 -281 500 -247
rect 590 -281 718 -247
<< metal1 >>
rect -804 419 804 425
rect -920 385 -874 397
rect -920 38 -914 385
rect -880 38 -874 385
rect -804 385 -792 419
rect 792 385 804 419
rect -804 379 804 385
rect -730 281 -578 287
rect -730 247 -718 281
rect -590 247 -578 281
rect -730 241 -578 247
rect -512 281 -360 287
rect -512 247 -500 281
rect -372 247 -360 281
rect -512 241 -360 247
rect -294 281 -142 287
rect -294 247 -282 281
rect -154 247 -142 281
rect -294 241 -142 247
rect -76 281 76 287
rect -76 247 -64 281
rect 64 247 76 281
rect -76 241 76 247
rect 142 281 294 287
rect 142 247 154 281
rect 282 247 294 281
rect 142 241 294 247
rect 360 281 512 287
rect 360 247 372 281
rect 500 247 512 281
rect 360 241 512 247
rect 578 281 730 287
rect 578 247 590 281
rect 718 247 730 281
rect 578 241 730 247
rect -920 26 -874 38
rect -786 171 -740 183
rect -786 21 -780 171
rect -746 21 -740 171
rect -786 9 -740 21
rect -350 171 -304 183
rect -350 21 -344 171
rect -310 21 -304 171
rect -350 9 -304 21
rect 86 171 132 183
rect 86 21 92 171
rect 126 21 132 171
rect 86 9 132 21
rect 522 171 568 183
rect 522 21 528 171
rect 562 21 568 171
rect 522 9 568 21
rect -568 -21 -522 -9
rect -568 -171 -562 -21
rect -528 -171 -522 -21
rect -568 -183 -522 -171
rect -132 -21 -86 -9
rect -132 -171 -126 -21
rect -92 -171 -86 -21
rect -132 -183 -86 -171
rect 304 -21 350 -9
rect 304 -171 310 -21
rect 344 -171 350 -21
rect 304 -183 350 -171
rect 740 -21 786 -9
rect 740 -171 746 -21
rect 780 -171 786 -21
rect 740 -183 786 -171
rect -730 -247 -578 -241
rect -730 -281 -718 -247
rect -590 -281 -578 -247
rect -730 -287 -578 -281
rect -512 -247 -360 -241
rect -512 -281 -500 -247
rect -372 -281 -360 -247
rect -512 -287 -360 -281
rect -294 -247 -142 -241
rect -294 -281 -282 -247
rect -154 -281 -142 -247
rect -294 -287 -142 -281
rect -76 -247 76 -241
rect -76 -281 -64 -247
rect 64 -281 76 -247
rect -76 -287 76 -281
rect 142 -247 294 -241
rect 142 -281 154 -247
rect 282 -281 294 -247
rect 142 -287 294 -281
rect 360 -247 512 -241
rect 360 -281 372 -247
rect 500 -281 512 -247
rect 360 -287 512 -281
rect 578 -247 730 -241
rect 578 -281 590 -247
rect 718 -281 730 -247
rect 578 -287 730 -281
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string FIXED_BBOX -897 -402 897 402
string parameters w 2.00 l 0.80 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl -45 viagr 0 viagt 90 viagb 0 viagate 100 viadrn -40 viasrc +40
string library sky130
<< end >>
