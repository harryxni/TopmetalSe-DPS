magic
tech sky130B
magscale 1 2
timestamp 1607712711
<< viali >>
rect 2911 1130 2945 1164
rect 2431 612 2465 646
<< metal1 >>
rect 0 4910 4992 4935
rect 0 4858 1544 4910
rect 1596 4858 1608 4910
rect 1660 4858 1672 4910
rect 1724 4858 1736 4910
rect 1788 4858 3211 4910
rect 3263 4858 3275 4910
rect 3327 4858 3339 4910
rect 3391 4858 3403 4910
rect 3455 4858 4992 4910
rect 0 4833 4992 4858
rect 0 3282 4992 3307
rect 0 3230 711 3282
rect 763 3230 775 3282
rect 827 3230 839 3282
rect 891 3230 903 3282
rect 955 3230 2378 3282
rect 2430 3230 2442 3282
rect 2494 3230 2506 3282
rect 2558 3230 2570 3282
rect 2622 3230 4044 3282
rect 4096 3230 4108 3282
rect 4160 3230 4172 3282
rect 4224 3230 4236 3282
rect 4288 3230 4992 3282
rect 0 3205 4992 3230
rect 0 1654 4992 1679
rect 0 1602 1544 1654
rect 1596 1602 1608 1654
rect 1660 1602 1672 1654
rect 1724 1602 1736 1654
rect 1788 1602 3211 1654
rect 3263 1602 3275 1654
rect 3327 1602 3339 1654
rect 3391 1602 3403 1654
rect 3455 1602 4992 1654
rect 0 1577 4992 1602
rect 592 1121 598 1173
rect 650 1161 656 1173
rect 2899 1164 2957 1170
rect 2899 1161 2911 1164
rect 650 1133 2911 1161
rect 650 1121 656 1133
rect 2899 1130 2911 1133
rect 2945 1130 2957 1164
rect 2899 1124 2957 1130
rect 2416 643 2422 655
rect 2377 615 2422 643
rect 2416 603 2422 615
rect 2474 603 2480 655
rect 0 26 4992 51
rect 0 -26 711 26
rect 763 -26 775 26
rect 827 -26 839 26
rect 891 -26 903 26
rect 955 -26 2378 26
rect 2430 -26 2442 26
rect 2494 -26 2506 26
rect 2558 -26 2570 26
rect 2622 -26 4044 26
rect 4096 -26 4108 26
rect 4160 -26 4172 26
rect 4224 -26 4236 26
rect 4288 -26 4992 26
rect 0 -51 4992 -26
<< via1 >>
rect 1544 4858 1596 4910
rect 1608 4858 1660 4910
rect 1672 4858 1724 4910
rect 1736 4858 1788 4910
rect 3211 4858 3263 4910
rect 3275 4858 3327 4910
rect 3339 4858 3391 4910
rect 3403 4858 3455 4910
rect 711 3230 763 3282
rect 775 3230 827 3282
rect 839 3230 891 3282
rect 903 3230 955 3282
rect 2378 3230 2430 3282
rect 2442 3230 2494 3282
rect 2506 3230 2558 3282
rect 2570 3230 2622 3282
rect 4044 3230 4096 3282
rect 4108 3230 4160 3282
rect 4172 3230 4224 3282
rect 4236 3230 4288 3282
rect 1544 1602 1596 1654
rect 1608 1602 1660 1654
rect 1672 1602 1724 1654
rect 1736 1602 1788 1654
rect 3211 1602 3263 1654
rect 3275 1602 3327 1654
rect 3339 1602 3391 1654
rect 3403 1602 3455 1654
rect 598 1121 650 1173
rect 2422 646 2474 655
rect 2422 612 2431 646
rect 2431 612 2465 646
rect 2465 612 2474 646
rect 2422 603 2474 612
rect 711 -26 763 26
rect 775 -26 827 26
rect 839 -26 891 26
rect 903 -26 955 26
rect 2378 -26 2430 26
rect 2442 -26 2494 26
rect 2506 -26 2558 26
rect 2570 -26 2622 26
rect 4044 -26 4096 26
rect 4108 -26 4160 26
rect 4172 -26 4224 26
rect 4236 -26 4288 26
<< metal2 >>
rect 1518 4912 1814 4935
rect 1574 4910 1598 4912
rect 1654 4910 1678 4912
rect 1734 4910 1758 4912
rect 1596 4858 1598 4910
rect 1660 4858 1672 4910
rect 1734 4858 1736 4910
rect 1574 4856 1598 4858
rect 1654 4856 1678 4858
rect 1734 4856 1758 4858
rect 1518 4833 1814 4856
rect 3185 4912 3481 4935
rect 3241 4910 3265 4912
rect 3321 4910 3345 4912
rect 3401 4910 3425 4912
rect 3263 4858 3265 4910
rect 3327 4858 3339 4910
rect 3401 4858 3403 4910
rect 3241 4856 3265 4858
rect 3321 4856 3345 4858
rect 3401 4856 3425 4858
rect 3185 4833 3481 4856
rect 4244 4200 4300 5000
rect 4258 3492 4286 4200
rect 4258 3464 4382 3492
rect 685 3284 981 3307
rect 741 3282 765 3284
rect 821 3282 845 3284
rect 901 3282 925 3284
rect 763 3230 765 3282
rect 827 3230 839 3282
rect 901 3230 903 3282
rect 741 3228 765 3230
rect 821 3228 845 3230
rect 901 3228 925 3230
rect 685 3205 981 3228
rect 2352 3284 2648 3307
rect 2408 3282 2432 3284
rect 2488 3282 2512 3284
rect 2568 3282 2592 3284
rect 2430 3230 2432 3282
rect 2494 3230 2506 3282
rect 2568 3230 2570 3282
rect 2408 3228 2432 3230
rect 2488 3228 2512 3230
rect 2568 3228 2592 3230
rect 2352 3205 2648 3228
rect 4018 3284 4314 3307
rect 4074 3282 4098 3284
rect 4154 3282 4178 3284
rect 4234 3282 4258 3284
rect 4096 3230 4098 3282
rect 4160 3230 4172 3282
rect 4234 3230 4236 3282
rect 4074 3228 4098 3230
rect 4154 3228 4178 3230
rect 4234 3228 4258 3230
rect 4018 3205 4314 3228
rect 1518 1656 1814 1679
rect 1574 1654 1598 1656
rect 1654 1654 1678 1656
rect 1734 1654 1758 1656
rect 1596 1602 1598 1654
rect 1660 1602 1672 1654
rect 1734 1602 1736 1654
rect 1574 1600 1598 1602
rect 1654 1600 1678 1602
rect 1734 1600 1758 1602
rect 1518 1577 1814 1600
rect 3185 1656 3481 1679
rect 3241 1654 3265 1656
rect 3321 1654 3345 1656
rect 3401 1654 3425 1656
rect 3263 1602 3265 1654
rect 3327 1602 3339 1654
rect 3401 1602 3403 1654
rect 3241 1600 3265 1602
rect 3321 1600 3345 1602
rect 3401 1600 3425 1602
rect 3185 1577 3481 1600
rect 598 1173 650 1179
rect 598 1115 650 1121
rect 610 800 638 1115
rect 596 0 652 800
rect 4354 703 4382 3464
rect 2420 694 2476 703
rect 2420 629 2422 638
rect 2474 629 2476 638
rect 4340 694 4396 703
rect 4340 629 4396 638
rect 2422 597 2474 603
rect 685 28 981 51
rect 741 26 765 28
rect 821 26 845 28
rect 901 26 925 28
rect 763 -26 765 26
rect 827 -26 839 26
rect 901 -26 903 26
rect 741 -28 765 -26
rect 821 -28 845 -26
rect 901 -28 925 -26
rect 685 -51 981 -28
rect 2352 28 2648 51
rect 2408 26 2432 28
rect 2488 26 2512 28
rect 2568 26 2592 28
rect 2430 -26 2432 26
rect 2494 -26 2506 26
rect 2568 -26 2570 26
rect 2408 -28 2432 -26
rect 2488 -28 2512 -26
rect 2568 -28 2592 -26
rect 2352 -51 2648 -28
rect 4018 28 4314 51
rect 4074 26 4098 28
rect 4154 26 4178 28
rect 4234 26 4258 28
rect 4096 -26 4098 26
rect 4160 -26 4172 26
rect 4234 -26 4236 26
rect 4074 -28 4098 -26
rect 4154 -28 4178 -26
rect 4234 -28 4258 -26
rect 4018 -51 4314 -28
<< via2 >>
rect 1518 4910 1574 4912
rect 1598 4910 1654 4912
rect 1678 4910 1734 4912
rect 1758 4910 1814 4912
rect 1518 4858 1544 4910
rect 1544 4858 1574 4910
rect 1598 4858 1608 4910
rect 1608 4858 1654 4910
rect 1678 4858 1724 4910
rect 1724 4858 1734 4910
rect 1758 4858 1788 4910
rect 1788 4858 1814 4910
rect 1518 4856 1574 4858
rect 1598 4856 1654 4858
rect 1678 4856 1734 4858
rect 1758 4856 1814 4858
rect 3185 4910 3241 4912
rect 3265 4910 3321 4912
rect 3345 4910 3401 4912
rect 3425 4910 3481 4912
rect 3185 4858 3211 4910
rect 3211 4858 3241 4910
rect 3265 4858 3275 4910
rect 3275 4858 3321 4910
rect 3345 4858 3391 4910
rect 3391 4858 3401 4910
rect 3425 4858 3455 4910
rect 3455 4858 3481 4910
rect 3185 4856 3241 4858
rect 3265 4856 3321 4858
rect 3345 4856 3401 4858
rect 3425 4856 3481 4858
rect 685 3282 741 3284
rect 765 3282 821 3284
rect 845 3282 901 3284
rect 925 3282 981 3284
rect 685 3230 711 3282
rect 711 3230 741 3282
rect 765 3230 775 3282
rect 775 3230 821 3282
rect 845 3230 891 3282
rect 891 3230 901 3282
rect 925 3230 955 3282
rect 955 3230 981 3282
rect 685 3228 741 3230
rect 765 3228 821 3230
rect 845 3228 901 3230
rect 925 3228 981 3230
rect 2352 3282 2408 3284
rect 2432 3282 2488 3284
rect 2512 3282 2568 3284
rect 2592 3282 2648 3284
rect 2352 3230 2378 3282
rect 2378 3230 2408 3282
rect 2432 3230 2442 3282
rect 2442 3230 2488 3282
rect 2512 3230 2558 3282
rect 2558 3230 2568 3282
rect 2592 3230 2622 3282
rect 2622 3230 2648 3282
rect 2352 3228 2408 3230
rect 2432 3228 2488 3230
rect 2512 3228 2568 3230
rect 2592 3228 2648 3230
rect 4018 3282 4074 3284
rect 4098 3282 4154 3284
rect 4178 3282 4234 3284
rect 4258 3282 4314 3284
rect 4018 3230 4044 3282
rect 4044 3230 4074 3282
rect 4098 3230 4108 3282
rect 4108 3230 4154 3282
rect 4178 3230 4224 3282
rect 4224 3230 4234 3282
rect 4258 3230 4288 3282
rect 4288 3230 4314 3282
rect 4018 3228 4074 3230
rect 4098 3228 4154 3230
rect 4178 3228 4234 3230
rect 4258 3228 4314 3230
rect 1518 1654 1574 1656
rect 1598 1654 1654 1656
rect 1678 1654 1734 1656
rect 1758 1654 1814 1656
rect 1518 1602 1544 1654
rect 1544 1602 1574 1654
rect 1598 1602 1608 1654
rect 1608 1602 1654 1654
rect 1678 1602 1724 1654
rect 1724 1602 1734 1654
rect 1758 1602 1788 1654
rect 1788 1602 1814 1654
rect 1518 1600 1574 1602
rect 1598 1600 1654 1602
rect 1678 1600 1734 1602
rect 1758 1600 1814 1602
rect 3185 1654 3241 1656
rect 3265 1654 3321 1656
rect 3345 1654 3401 1656
rect 3425 1654 3481 1656
rect 3185 1602 3211 1654
rect 3211 1602 3241 1654
rect 3265 1602 3275 1654
rect 3275 1602 3321 1654
rect 3345 1602 3391 1654
rect 3391 1602 3401 1654
rect 3425 1602 3455 1654
rect 3455 1602 3481 1654
rect 3185 1600 3241 1602
rect 3265 1600 3321 1602
rect 3345 1600 3401 1602
rect 3425 1600 3481 1602
rect 2420 655 2476 694
rect 2420 638 2422 655
rect 2422 638 2474 655
rect 2474 638 2476 655
rect 4340 638 4396 694
rect 685 26 741 28
rect 765 26 821 28
rect 845 26 901 28
rect 925 26 981 28
rect 685 -26 711 26
rect 711 -26 741 26
rect 765 -26 775 26
rect 775 -26 821 26
rect 845 -26 891 26
rect 891 -26 901 26
rect 925 -26 955 26
rect 955 -26 981 26
rect 685 -28 741 -26
rect 765 -28 821 -26
rect 845 -28 901 -26
rect 925 -28 981 -26
rect 2352 26 2408 28
rect 2432 26 2488 28
rect 2512 26 2568 28
rect 2592 26 2648 28
rect 2352 -26 2378 26
rect 2378 -26 2408 26
rect 2432 -26 2442 26
rect 2442 -26 2488 26
rect 2512 -26 2558 26
rect 2558 -26 2568 26
rect 2592 -26 2622 26
rect 2622 -26 2648 26
rect 2352 -28 2408 -26
rect 2432 -28 2488 -26
rect 2512 -28 2568 -26
rect 2592 -28 2648 -26
rect 4018 26 4074 28
rect 4098 26 4154 28
rect 4178 26 4234 28
rect 4258 26 4314 28
rect 4018 -26 4044 26
rect 4044 -26 4074 26
rect 4098 -26 4108 26
rect 4108 -26 4154 26
rect 4178 -26 4224 26
rect 4224 -26 4234 26
rect 4258 -26 4288 26
rect 4288 -26 4314 26
rect 4018 -28 4074 -26
rect 4098 -28 4154 -26
rect 4178 -28 4234 -26
rect 4258 -28 4314 -26
<< metal3 >>
rect 1506 4916 1826 4917
rect 1506 4852 1514 4916
rect 1578 4852 1594 4916
rect 1658 4852 1674 4916
rect 1738 4852 1754 4916
rect 1818 4852 1826 4916
rect 1506 4851 1826 4852
rect 3173 4916 3493 4917
rect 3173 4852 3181 4916
rect 3245 4852 3261 4916
rect 3325 4852 3341 4916
rect 3405 4852 3421 4916
rect 3485 4852 3493 4916
rect 3173 4851 3493 4852
rect 673 3288 993 3289
rect 673 3224 681 3288
rect 745 3224 761 3288
rect 825 3224 841 3288
rect 905 3224 921 3288
rect 985 3224 993 3288
rect 673 3223 993 3224
rect 2340 3288 2660 3289
rect 2340 3224 2348 3288
rect 2412 3224 2428 3288
rect 2492 3224 2508 3288
rect 2572 3224 2588 3288
rect 2652 3224 2660 3288
rect 2340 3223 2660 3224
rect 4006 3288 4326 3289
rect 4006 3224 4014 3288
rect 4078 3224 4094 3288
rect 4158 3224 4174 3288
rect 4238 3224 4254 3288
rect 4318 3224 4326 3288
rect 4006 3223 4326 3224
rect 1506 1660 1826 1661
rect 1506 1596 1514 1660
rect 1578 1596 1594 1660
rect 1658 1596 1674 1660
rect 1738 1596 1754 1660
rect 1818 1596 1826 1660
rect 1506 1595 1826 1596
rect 3173 1660 3493 1661
rect 3173 1596 3181 1660
rect 3245 1596 3261 1660
rect 3325 1596 3341 1660
rect 3405 1596 3421 1660
rect 3485 1596 3493 1660
rect 3173 1595 3493 1596
rect 2415 696 2481 699
rect 4335 696 4401 699
rect 2415 694 4401 696
rect 2415 638 2420 694
rect 2476 638 4340 694
rect 4396 638 4401 694
rect 2415 636 4401 638
rect 2415 633 2481 636
rect 4335 633 4401 636
rect 673 32 993 33
rect 673 -32 681 32
rect 745 -32 761 32
rect 825 -32 841 32
rect 905 -32 921 32
rect 985 -32 993 32
rect 673 -33 993 -32
rect 2340 32 2660 33
rect 2340 -32 2348 32
rect 2412 -32 2428 32
rect 2492 -32 2508 32
rect 2572 -32 2588 32
rect 2652 -32 2660 32
rect 2340 -33 2660 -32
rect 4006 32 4326 33
rect 4006 -32 4014 32
rect 4078 -32 4094 32
rect 4158 -32 4174 32
rect 4238 -32 4254 32
rect 4318 -32 4326 32
rect 4006 -33 4326 -32
<< via3 >>
rect 1514 4912 1578 4916
rect 1514 4856 1518 4912
rect 1518 4856 1574 4912
rect 1574 4856 1578 4912
rect 1514 4852 1578 4856
rect 1594 4912 1658 4916
rect 1594 4856 1598 4912
rect 1598 4856 1654 4912
rect 1654 4856 1658 4912
rect 1594 4852 1658 4856
rect 1674 4912 1738 4916
rect 1674 4856 1678 4912
rect 1678 4856 1734 4912
rect 1734 4856 1738 4912
rect 1674 4852 1738 4856
rect 1754 4912 1818 4916
rect 1754 4856 1758 4912
rect 1758 4856 1814 4912
rect 1814 4856 1818 4912
rect 1754 4852 1818 4856
rect 3181 4912 3245 4916
rect 3181 4856 3185 4912
rect 3185 4856 3241 4912
rect 3241 4856 3245 4912
rect 3181 4852 3245 4856
rect 3261 4912 3325 4916
rect 3261 4856 3265 4912
rect 3265 4856 3321 4912
rect 3321 4856 3325 4912
rect 3261 4852 3325 4856
rect 3341 4912 3405 4916
rect 3341 4856 3345 4912
rect 3345 4856 3401 4912
rect 3401 4856 3405 4912
rect 3341 4852 3405 4856
rect 3421 4912 3485 4916
rect 3421 4856 3425 4912
rect 3425 4856 3481 4912
rect 3481 4856 3485 4912
rect 3421 4852 3485 4856
rect 681 3284 745 3288
rect 681 3228 685 3284
rect 685 3228 741 3284
rect 741 3228 745 3284
rect 681 3224 745 3228
rect 761 3284 825 3288
rect 761 3228 765 3284
rect 765 3228 821 3284
rect 821 3228 825 3284
rect 761 3224 825 3228
rect 841 3284 905 3288
rect 841 3228 845 3284
rect 845 3228 901 3284
rect 901 3228 905 3284
rect 841 3224 905 3228
rect 921 3284 985 3288
rect 921 3228 925 3284
rect 925 3228 981 3284
rect 981 3228 985 3284
rect 921 3224 985 3228
rect 2348 3284 2412 3288
rect 2348 3228 2352 3284
rect 2352 3228 2408 3284
rect 2408 3228 2412 3284
rect 2348 3224 2412 3228
rect 2428 3284 2492 3288
rect 2428 3228 2432 3284
rect 2432 3228 2488 3284
rect 2488 3228 2492 3284
rect 2428 3224 2492 3228
rect 2508 3284 2572 3288
rect 2508 3228 2512 3284
rect 2512 3228 2568 3284
rect 2568 3228 2572 3284
rect 2508 3224 2572 3228
rect 2588 3284 2652 3288
rect 2588 3228 2592 3284
rect 2592 3228 2648 3284
rect 2648 3228 2652 3284
rect 2588 3224 2652 3228
rect 4014 3284 4078 3288
rect 4014 3228 4018 3284
rect 4018 3228 4074 3284
rect 4074 3228 4078 3284
rect 4014 3224 4078 3228
rect 4094 3284 4158 3288
rect 4094 3228 4098 3284
rect 4098 3228 4154 3284
rect 4154 3228 4158 3284
rect 4094 3224 4158 3228
rect 4174 3284 4238 3288
rect 4174 3228 4178 3284
rect 4178 3228 4234 3284
rect 4234 3228 4238 3284
rect 4174 3224 4238 3228
rect 4254 3284 4318 3288
rect 4254 3228 4258 3284
rect 4258 3228 4314 3284
rect 4314 3228 4318 3284
rect 4254 3224 4318 3228
rect 1514 1656 1578 1660
rect 1514 1600 1518 1656
rect 1518 1600 1574 1656
rect 1574 1600 1578 1656
rect 1514 1596 1578 1600
rect 1594 1656 1658 1660
rect 1594 1600 1598 1656
rect 1598 1600 1654 1656
rect 1654 1600 1658 1656
rect 1594 1596 1658 1600
rect 1674 1656 1738 1660
rect 1674 1600 1678 1656
rect 1678 1600 1734 1656
rect 1734 1600 1738 1656
rect 1674 1596 1738 1600
rect 1754 1656 1818 1660
rect 1754 1600 1758 1656
rect 1758 1600 1814 1656
rect 1814 1600 1818 1656
rect 1754 1596 1818 1600
rect 3181 1656 3245 1660
rect 3181 1600 3185 1656
rect 3185 1600 3241 1656
rect 3241 1600 3245 1656
rect 3181 1596 3245 1600
rect 3261 1656 3325 1660
rect 3261 1600 3265 1656
rect 3265 1600 3321 1656
rect 3321 1600 3325 1656
rect 3261 1596 3325 1600
rect 3341 1656 3405 1660
rect 3341 1600 3345 1656
rect 3345 1600 3401 1656
rect 3401 1600 3405 1656
rect 3341 1596 3405 1600
rect 3421 1656 3485 1660
rect 3421 1600 3425 1656
rect 3425 1600 3481 1656
rect 3481 1600 3485 1656
rect 3421 1596 3485 1600
rect 681 28 745 32
rect 681 -28 685 28
rect 685 -28 741 28
rect 741 -28 745 28
rect 681 -32 745 -28
rect 761 28 825 32
rect 761 -28 765 28
rect 765 -28 821 28
rect 821 -28 825 28
rect 761 -32 825 -28
rect 841 28 905 32
rect 841 -28 845 28
rect 845 -28 901 28
rect 901 -28 905 28
rect 841 -32 905 -28
rect 921 28 985 32
rect 921 -28 925 28
rect 925 -28 981 28
rect 981 -28 985 28
rect 921 -32 985 -28
rect 2348 28 2412 32
rect 2348 -28 2352 28
rect 2352 -28 2408 28
rect 2408 -28 2412 28
rect 2348 -32 2412 -28
rect 2428 28 2492 32
rect 2428 -28 2432 28
rect 2432 -28 2488 28
rect 2488 -28 2492 28
rect 2428 -32 2492 -28
rect 2508 28 2572 32
rect 2508 -28 2512 28
rect 2512 -28 2568 28
rect 2568 -28 2572 28
rect 2508 -32 2572 -28
rect 2588 28 2652 32
rect 2588 -28 2592 28
rect 2592 -28 2648 28
rect 2648 -28 2652 28
rect 2588 -32 2652 -28
rect 4014 28 4078 32
rect 4014 -28 4018 28
rect 4018 -28 4074 28
rect 4074 -28 4078 28
rect 4014 -32 4078 -28
rect 4094 28 4158 32
rect 4094 -28 4098 28
rect 4098 -28 4154 28
rect 4154 -28 4158 28
rect 4094 -32 4158 -28
rect 4174 28 4238 32
rect 4174 -28 4178 28
rect 4178 -28 4234 28
rect 4234 -28 4238 28
rect 4174 -32 4238 -28
rect 4254 28 4318 32
rect 4254 -28 4258 28
rect 4258 -28 4314 28
rect 4314 -28 4318 28
rect 4254 -32 4318 -28
<< metal4 >>
rect 673 4233 993 4935
rect 673 3997 715 4233
rect 951 3997 993 4233
rect 673 3288 993 3997
rect 673 3224 681 3288
rect 745 3224 761 3288
rect 825 3224 841 3288
rect 905 3224 921 3288
rect 985 3224 993 3288
rect 673 2567 993 3224
rect 673 2331 715 2567
rect 951 2331 993 2567
rect 673 900 993 2331
rect 673 664 715 900
rect 951 664 993 900
rect 673 32 993 664
rect 673 -32 681 32
rect 745 -32 761 32
rect 825 -32 841 32
rect 905 -32 921 32
rect 985 -32 993 32
rect 673 -51 993 -32
rect 1506 4916 1827 4935
rect 1506 4852 1514 4916
rect 1578 4852 1594 4916
rect 1658 4852 1674 4916
rect 1738 4852 1754 4916
rect 1818 4852 1827 4916
rect 1506 3400 1827 4852
rect 1506 3164 1548 3400
rect 1784 3164 1827 3400
rect 1506 1733 1827 3164
rect 1506 1660 1548 1733
rect 1784 1660 1827 1733
rect 1506 1596 1514 1660
rect 1818 1596 1827 1660
rect 1506 1497 1548 1596
rect 1784 1497 1827 1596
rect 1506 -51 1827 1497
rect 2340 4233 2660 4935
rect 2340 3997 2382 4233
rect 2618 3997 2660 4233
rect 2340 3288 2660 3997
rect 2340 3224 2348 3288
rect 2412 3224 2428 3288
rect 2492 3224 2508 3288
rect 2572 3224 2588 3288
rect 2652 3224 2660 3288
rect 2340 2567 2660 3224
rect 2340 2331 2382 2567
rect 2618 2331 2660 2567
rect 2340 900 2660 2331
rect 2340 664 2382 900
rect 2618 664 2660 900
rect 2340 32 2660 664
rect 2340 -32 2348 32
rect 2412 -32 2428 32
rect 2492 -32 2508 32
rect 2572 -32 2588 32
rect 2652 -32 2660 32
rect 2340 -51 2660 -32
rect 3173 4916 3493 4935
rect 3173 4852 3181 4916
rect 3245 4852 3261 4916
rect 3325 4852 3341 4916
rect 3405 4852 3421 4916
rect 3485 4852 3493 4916
rect 3173 3400 3493 4852
rect 3173 3164 3215 3400
rect 3451 3164 3493 3400
rect 3173 1733 3493 3164
rect 3173 1660 3215 1733
rect 3451 1660 3493 1733
rect 3173 1596 3181 1660
rect 3485 1596 3493 1660
rect 3173 1497 3215 1596
rect 3451 1497 3493 1596
rect 3173 -51 3493 1497
rect 4006 4233 4327 4935
rect 4006 3997 4048 4233
rect 4284 3997 4327 4233
rect 4006 3288 4327 3997
rect 4006 3224 4014 3288
rect 4078 3224 4094 3288
rect 4158 3224 4174 3288
rect 4238 3224 4254 3288
rect 4318 3224 4327 3288
rect 4006 2567 4327 3224
rect 4006 2331 4048 2567
rect 4284 2331 4327 2567
rect 4006 900 4327 2331
rect 4006 664 4048 900
rect 4284 664 4327 900
rect 4006 32 4327 664
rect 4006 -32 4014 32
rect 4078 -32 4094 32
rect 4158 -32 4174 32
rect 4238 -32 4254 32
rect 4318 -32 4327 32
rect 4006 -51 4327 -32
<< via4 >>
rect 715 3997 951 4233
rect 715 2331 951 2567
rect 715 664 951 900
rect 1548 3164 1784 3400
rect 1548 1660 1784 1733
rect 1548 1596 1578 1660
rect 1578 1596 1594 1660
rect 1594 1596 1658 1660
rect 1658 1596 1674 1660
rect 1674 1596 1738 1660
rect 1738 1596 1754 1660
rect 1754 1596 1784 1660
rect 1548 1497 1784 1596
rect 2382 3997 2618 4233
rect 2382 2331 2618 2567
rect 2382 664 2618 900
rect 3215 3164 3451 3400
rect 3215 1660 3451 1733
rect 3215 1596 3245 1660
rect 3245 1596 3261 1660
rect 3261 1596 3325 1660
rect 3325 1596 3341 1660
rect 3341 1596 3405 1660
rect 3405 1596 3421 1660
rect 3421 1596 3451 1660
rect 3215 1497 3451 1596
rect 4048 3997 4284 4233
rect 4048 2331 4284 2567
rect 4048 664 4284 900
<< metal5 >>
rect 0 4233 4992 4276
rect 0 3997 715 4233
rect 951 3997 2382 4233
rect 2618 3997 4048 4233
rect 4284 3997 4992 4233
rect 0 3955 4992 3997
rect 0 3400 4992 3442
rect 0 3164 1548 3400
rect 1784 3164 3215 3400
rect 3451 3164 4992 3400
rect 0 3122 4992 3164
rect 0 2567 4992 2609
rect 0 2331 715 2567
rect 951 2331 2382 2567
rect 2618 2331 4048 2567
rect 4284 2331 4992 2567
rect 0 2289 4992 2331
rect 0 1733 4992 1776
rect 0 1497 1548 1733
rect 1784 1497 3215 1733
rect 3451 1497 4992 1733
rect 0 1455 4992 1497
rect 0 900 4992 942
rect 0 664 715 900
rect 951 664 2382 900
rect 2618 664 4048 900
rect 4284 664 4992 900
rect 0 622 4992 664
use sky130_fd_sc_hvl__decap_8  FILLER_0_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1607116011
transform 1 0 0 0 -1 814
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_8
timestamp 1607116011
transform 1 0 768 0 -1 814
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_0_16 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1607116011
transform 1 0 1536 0 -1 814
box -66 -23 450 897
use sky130_fd_sc_hvl__lsbufhv2lv_1  lvlshiftdown $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1607116011
transform 1 0 2208 0 -1 1628
box -66 -23 1698 1651
use sky130_fd_sc_hvl__fill_2  FILLER_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1607116011
transform 1 0 1920 0 -1 814
box -66 -23 258 897
use sky130_fd_sc_hvl__fill_1  FILLER_0_22 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1607116011
transform 1 0 2112 0 -1 814
box -66 -23 162 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_40
timestamp 1607116011
transform 1 0 3840 0 -1 814
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_0_48
timestamp 1607116011
transform 1 0 4608 0 -1 814
box -66 -23 450 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_0
timestamp 1607116011
transform 1 0 0 0 1 1628
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_8
timestamp 1607116011
transform 1 0 768 0 1 1628
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_16
timestamp 1607116011
transform 1 0 1536 0 1 1628
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_0
timestamp 1607116011
transform 1 0 0 0 -1 4070
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_8
timestamp 1607116011
transform 1 0 768 0 -1 4070
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_16
timestamp 1607116011
transform 1 0 1536 0 -1 4070
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_24
timestamp 1607116011
transform 1 0 2304 0 1 1628
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_32
timestamp 1607116011
transform 1 0 3072 0 1 1628
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_24
timestamp 1607116011
transform 1 0 2304 0 -1 4070
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_32
timestamp 1607116011
transform 1 0 3072 0 -1 4070
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_40
timestamp 1607116011
transform 1 0 3840 0 1 1628
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_1_48
timestamp 1607116011
transform 1 0 4608 0 1 1628
box -66 -23 450 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_40
timestamp 1607116011
transform 1 0 3840 0 -1 4070
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_2_48
timestamp 1607116011
transform 1 0 4608 0 -1 4070
box -66 -23 450 897
<< labels >>
rlabel metal2 s 4244 4200 4300 5000 6 A
port 0 nsew signal input
rlabel metal2 s 596 0 652 800 6 X
port 1 nsew signal tristate
rlabel metal4 s 4007 -51 4327 4935 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 2340 -51 2660 4935 6 VPWR
port 3 nsew power bidirectional
rlabel metal4 s 673 -51 993 4935 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 3956 4992 4276 6 VPWR
port 5 nsew power bidirectional
rlabel metal5 s 0 2289 4992 2609 6 VPWR
port 6 nsew power bidirectional
rlabel metal5 s 0 622 4992 942 6 VPWR
port 7 nsew power bidirectional
rlabel metal4 s 3173 -51 3493 4935 6 VGND
port 8 nsew ground bidirectional
rlabel metal4 s 1507 -51 1827 4935 6 VGND
port 9 nsew ground bidirectional
rlabel metal5 s 0 3122 4992 3442 6 VGND
port 10 nsew ground bidirectional
rlabel metal5 s 0 1456 4992 1776 6 VGND
port 11 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 5000 5000
<< end >>
