magic
tech sky130B
magscale 1 2
timestamp 1661984010
<< nwell >>
rect 1010 -1030 1930 -510
<< nmos >>
rect 7150 -600 8150 -400
rect 8350 -600 9350 -400
rect 9480 -600 10480 -400
rect 8460 -1450 8544 -1250
rect 9580 -1450 9680 -1250
<< pmoslvt >>
rect 1280 -960 1480 -760
<< nmoslvt >>
rect 2360 -1410 2560 -1170
rect 2870 -1410 3070 -1170
rect 3230 -1330 4830 -930
rect 5230 -1330 6830 -930
rect 7630 -1420 7830 -1220
<< ndiff >>
rect 7150 -320 8150 -300
rect 7150 -380 7170 -320
rect 8130 -380 8150 -320
rect 7150 -400 8150 -380
rect 8350 -320 9350 -300
rect 8350 -380 8370 -320
rect 9330 -380 9350 -320
rect 8350 -400 9350 -380
rect 9480 -320 10480 -300
rect 9480 -380 9500 -320
rect 10460 -380 10480 -320
rect 9480 -400 10480 -380
rect 7150 -640 8150 -600
rect 7150 -700 7270 -640
rect 3230 -810 4830 -790
rect 3230 -910 3250 -810
rect 4810 -910 4830 -810
rect 3230 -930 4830 -910
rect 5230 -810 6830 -790
rect 5230 -910 5250 -810
rect 6810 -910 6830 -810
rect 7220 -810 7270 -700
rect 8100 -810 8150 -640
rect 8350 -640 9350 -600
rect 8350 -700 8470 -640
rect 7220 -830 8150 -810
rect 8420 -810 8470 -700
rect 9300 -810 9350 -640
rect 9480 -640 10480 -600
rect 9480 -700 9600 -640
rect 8420 -830 9350 -810
rect 9550 -810 9600 -700
rect 10430 -810 10480 -640
rect 9550 -830 10480 -810
rect 5230 -930 6830 -910
rect 2360 -1110 2560 -1100
rect 2360 -1150 2380 -1110
rect 2540 -1150 2560 -1110
rect 2360 -1170 2560 -1150
rect 2870 -1110 3070 -1100
rect 2870 -1150 2890 -1110
rect 3050 -1150 3070 -1110
rect 2870 -1170 3070 -1150
rect 8460 -1060 8544 -1050
rect 7630 -1140 7830 -1130
rect 7630 -1200 7650 -1140
rect 7810 -1200 7830 -1140
rect 7630 -1220 7830 -1200
rect 3230 -1350 4830 -1330
rect 2360 -1430 2560 -1410
rect 2360 -1470 2380 -1430
rect 2540 -1470 2560 -1430
rect 2360 -1480 2560 -1470
rect 2870 -1430 3070 -1410
rect 2870 -1470 2890 -1430
rect 3050 -1470 3070 -1430
rect 3230 -1450 3250 -1350
rect 4810 -1450 4830 -1350
rect 3230 -1460 4830 -1450
rect 5230 -1350 6830 -1330
rect 5230 -1450 5250 -1350
rect 6810 -1450 6830 -1350
rect 8460 -1230 8480 -1060
rect 8530 -1230 8544 -1060
rect 9590 -1060 9674 -1050
rect 9590 -1130 9610 -1060
rect 8460 -1250 8544 -1230
rect 9580 -1230 9610 -1130
rect 9660 -1130 9674 -1060
rect 9660 -1230 9680 -1130
rect 9580 -1250 9680 -1230
rect 5230 -1460 6830 -1450
rect 2870 -1480 3070 -1470
rect 7630 -1440 7830 -1420
rect 7630 -1530 7650 -1440
rect 7810 -1530 7830 -1440
rect 7630 -1590 7830 -1530
rect 8460 -1470 8544 -1450
rect 8460 -1640 8480 -1470
rect 8530 -1640 8544 -1470
rect 9580 -1470 9680 -1450
rect 9580 -1580 9600 -1470
rect 9660 -1580 9680 -1470
rect 9580 -1590 9680 -1580
rect 8460 -1650 8544 -1640
<< pdiff >>
rect 1190 -780 1280 -760
rect 1190 -940 1200 -780
rect 1260 -940 1280 -780
rect 1190 -960 1280 -940
rect 1480 -780 1590 -760
rect 1480 -940 1500 -780
rect 1560 -940 1590 -780
rect 1480 -960 1590 -940
<< ndiffc >>
rect 7170 -380 8130 -320
rect 8370 -380 9330 -320
rect 9500 -380 10460 -320
rect 3250 -910 4810 -810
rect 5250 -910 6810 -810
rect 7270 -810 8100 -640
rect 8470 -810 9300 -640
rect 9600 -810 10430 -640
rect 2380 -1150 2540 -1110
rect 2890 -1150 3050 -1110
rect 7650 -1200 7810 -1140
rect 2380 -1470 2540 -1430
rect 2890 -1470 3050 -1430
rect 3250 -1450 4810 -1350
rect 5250 -1450 6810 -1350
rect 8480 -1230 8530 -1060
rect 9610 -1230 9660 -1060
rect 7650 -1530 7810 -1440
rect 8480 -1640 8530 -1470
rect 9600 -1580 9660 -1470
<< pdiffc >>
rect 1200 -940 1260 -780
rect 1500 -940 1560 -780
<< psubdiff >>
rect 5230 -1490 6830 -1460
rect 5230 -1580 5260 -1490
rect 6800 -1580 6830 -1490
rect 5230 -1600 6830 -1580
<< nsubdiff >>
rect 1090 -790 1190 -760
rect 1090 -930 1110 -790
rect 1160 -930 1190 -790
rect 1090 -960 1190 -930
<< psubdiffcont >>
rect 5260 -1580 6800 -1490
<< nsubdiffcont >>
rect 1110 -930 1160 -790
<< poly >>
rect 10620 -400 10850 -380
rect 7120 -600 7150 -400
rect 8150 -600 8350 -400
rect 9350 -600 9480 -400
rect 10480 -410 10850 -400
rect 10480 -590 10640 -410
rect 10820 -590 10850 -410
rect 10480 -600 10850 -590
rect 1280 -760 1480 -730
rect 10620 -620 10850 -600
rect 1280 -990 1480 -960
rect 1280 -1050 1360 -990
rect 1280 -1110 1290 -1050
rect 1350 -1110 1360 -1050
rect 1280 -1130 1360 -1110
rect 2330 -1330 2360 -1170
rect 2230 -1340 2360 -1330
rect 2230 -1400 2250 -1340
rect 2310 -1400 2360 -1340
rect 2230 -1410 2360 -1400
rect 2560 -1410 2590 -1170
rect 2840 -1330 2870 -1170
rect 2740 -1340 2870 -1330
rect 2740 -1400 2760 -1340
rect 2820 -1400 2870 -1340
rect 2740 -1410 2870 -1400
rect 3070 -1410 3100 -1170
rect 3200 -1330 3230 -930
rect 4830 -1180 4860 -930
rect 4830 -1200 5020 -1180
rect 4830 -1310 4890 -1200
rect 5000 -1310 5020 -1200
rect 4830 -1330 5020 -1310
rect 5200 -1330 5230 -930
rect 6830 -1180 6860 -930
rect 6830 -1200 7020 -1180
rect 6830 -1310 6890 -1200
rect 7000 -1310 7020 -1200
rect 6830 -1330 7020 -1310
rect 7600 -1420 7630 -1220
rect 7830 -1300 7860 -1220
rect 7830 -1310 8011 -1300
rect 7830 -1360 7945 -1310
rect 7995 -1360 8011 -1310
rect 7830 -1370 8011 -1360
rect 7830 -1420 7860 -1370
rect 8430 -1450 8460 -1250
rect 8544 -1330 8570 -1250
rect 8630 -1330 8710 -1324
rect 8544 -1340 8710 -1330
rect 8544 -1400 8640 -1340
rect 8700 -1400 8710 -1340
rect 8544 -1410 8710 -1400
rect 8544 -1450 8570 -1410
rect 8630 -1416 8710 -1410
rect 9550 -1450 9580 -1250
rect 9680 -1330 9710 -1250
rect 9760 -1330 9840 -1324
rect 9680 -1340 9840 -1330
rect 9680 -1400 9770 -1340
rect 9830 -1400 9840 -1340
rect 9680 -1410 9840 -1400
rect 9680 -1450 9710 -1410
rect 9760 -1416 9840 -1410
<< polycont >>
rect 10640 -590 10820 -410
rect 1290 -1110 1350 -1050
rect 2250 -1400 2310 -1340
rect 2760 -1400 2820 -1340
rect 4890 -1310 5000 -1200
rect 6890 -1310 7000 -1200
rect 7945 -1360 7995 -1310
rect 8640 -1400 8700 -1340
rect 9770 -1400 9830 -1340
<< locali >>
rect 7150 -200 8150 -180
rect 7150 -380 7170 -200
rect 8130 -380 8150 -200
rect 8350 -200 9350 -180
rect 8350 -380 8370 -200
rect 9330 -380 9350 -200
rect 9480 -200 10480 -180
rect 9480 -380 9500 -200
rect 10460 -380 10480 -200
rect 10620 -400 10850 -380
rect 10620 -600 10630 -400
rect 10830 -600 10850 -400
rect 10620 -620 10850 -600
rect 7250 -640 8120 -620
rect 1090 -770 1190 -740
rect 1090 -780 1280 -770
rect 1090 -790 1200 -780
rect 1090 -930 1110 -790
rect 1160 -930 1200 -790
rect 1090 -940 1200 -930
rect 1260 -940 1280 -780
rect 1090 -950 1280 -940
rect 1480 -780 1580 -770
rect 1480 -940 1500 -780
rect 1560 -940 1580 -780
rect 3230 -810 5150 -790
rect 3230 -910 3250 -810
rect 4810 -910 5150 -810
rect 5230 -810 7150 -790
rect 5230 -910 5250 -810
rect 6810 -910 7150 -810
rect 1480 -950 1580 -940
rect 1500 -1040 1580 -950
rect 1090 -1050 1580 -1040
rect 1090 -1120 1110 -1050
rect 1200 -1110 1290 -1050
rect 1350 -1110 1470 -1050
rect 1200 -1120 1470 -1110
rect 1090 -1130 1580 -1120
rect 2250 -1150 2380 -1090
rect 2540 -1150 2560 -1090
rect 2760 -1150 2890 -1090
rect 3050 -1150 3070 -1090
rect 2250 -1330 2310 -1150
rect 2760 -1330 2820 -1150
rect 5040 -1200 5150 -910
rect 7040 -1200 7150 -910
rect 7250 -910 7270 -640
rect 8100 -910 8120 -640
rect 7250 -920 8120 -910
rect 8450 -640 9320 -620
rect 8450 -910 8470 -640
rect 9300 -910 9320 -640
rect 8450 -920 9320 -910
rect 9580 -640 10450 -620
rect 9580 -910 9600 -640
rect 10430 -910 10450 -640
rect 9580 -920 10450 -910
rect 7630 -1200 7650 -1000
rect 7810 -1055 7830 -1000
rect 8450 -1050 8560 -1030
rect 7810 -1125 8005 -1055
rect 7810 -1200 7830 -1125
rect 4860 -1310 4890 -1200
rect 5000 -1210 5150 -1200
rect 5120 -1300 5150 -1210
rect 5000 -1310 5150 -1300
rect 6860 -1310 6890 -1200
rect 7000 -1210 7150 -1200
rect 7120 -1300 7150 -1210
rect 7000 -1310 7150 -1300
rect 7935 -1215 8005 -1125
rect 8450 -1210 8460 -1050
rect 8550 -1140 8560 -1050
rect 9580 -1050 9690 -1030
rect 8550 -1210 8710 -1140
rect 8450 -1230 8480 -1210
rect 8530 -1220 8710 -1210
rect 8530 -1230 8560 -1220
rect 7935 -1310 8005 -1285
rect 2180 -1340 2310 -1330
rect 2220 -1400 2250 -1340
rect 2180 -1410 2310 -1400
rect 2600 -1340 2820 -1330
rect 2600 -1400 2620 -1340
rect 2730 -1400 2760 -1340
rect 2600 -1410 2820 -1400
rect 3230 -1350 4820 -1330
rect 2250 -1420 2310 -1410
rect 2360 -1430 2560 -1410
rect 2760 -1420 2820 -1410
rect 2360 -1470 2380 -1430
rect 2540 -1470 2560 -1430
rect 2360 -1550 2560 -1470
rect 2360 -1580 2370 -1550
rect 2550 -1580 2560 -1550
rect 2870 -1430 3070 -1410
rect 2870 -1470 2890 -1430
rect 3050 -1470 3070 -1430
rect 2870 -1550 3070 -1470
rect 2870 -1580 2880 -1550
rect 3060 -1580 3070 -1550
rect 3230 -1450 3250 -1350
rect 4810 -1450 4820 -1350
rect 3230 -1460 4820 -1450
rect 5230 -1350 6820 -1330
rect 5230 -1450 5250 -1350
rect 6810 -1450 6820 -1350
rect 7935 -1360 7945 -1310
rect 7995 -1360 8005 -1310
rect 8630 -1240 8710 -1220
rect 9580 -1210 9590 -1050
rect 9680 -1140 9690 -1050
rect 9680 -1210 9840 -1140
rect 9580 -1230 9610 -1210
rect 9660 -1220 9840 -1210
rect 9660 -1230 9690 -1220
rect 8630 -1340 8710 -1320
rect 9760 -1240 9840 -1220
rect 9760 -1340 9840 -1320
rect 7935 -1370 8005 -1360
rect 7945 -1376 7995 -1370
rect 8624 -1400 8640 -1340
rect 8700 -1400 8716 -1340
rect 9754 -1400 9770 -1340
rect 9830 -1400 9846 -1340
rect 8630 -1410 8710 -1400
rect 9760 -1410 9840 -1400
rect 3230 -1550 4830 -1460
rect 3230 -1580 3250 -1550
rect 4810 -1580 4830 -1550
rect 5230 -1476 6820 -1450
rect 5230 -1490 6830 -1476
rect 5230 -1540 5260 -1490
rect 6800 -1540 6830 -1490
rect 5230 -1580 5250 -1540
rect 6810 -1580 6830 -1540
rect 7630 -1530 7650 -1440
rect 7810 -1530 7830 -1440
rect 7630 -1580 7830 -1530
rect 8460 -1470 8544 -1450
rect 8460 -1580 8480 -1470
rect 8530 -1580 8544 -1470
rect 9580 -1470 9680 -1450
rect 9580 -1580 9600 -1470
rect 9660 -1580 9680 -1470
<< viali >>
rect 880 -710 1910 -240
rect 7170 -320 8130 -200
rect 7170 -370 8130 -320
rect 8370 -320 9330 -200
rect 8370 -370 9330 -320
rect 9500 -320 10460 -200
rect 9500 -370 10460 -320
rect 10630 -410 10830 -400
rect 10630 -590 10640 -410
rect 10640 -590 10820 -410
rect 10820 -590 10830 -410
rect 10630 -600 10830 -590
rect 1090 -740 1190 -710
rect 3250 -900 4810 -810
rect 5250 -900 6810 -810
rect 1110 -1120 1200 -1050
rect 1470 -1120 1580 -1050
rect 2380 -1110 2540 -1090
rect 2380 -1130 2540 -1110
rect 2890 -1110 3050 -1090
rect 2890 -1140 3050 -1110
rect 7270 -810 8100 -640
rect 7270 -910 8100 -810
rect 8470 -810 9300 -640
rect 8470 -910 9300 -810
rect 9600 -810 10430 -640
rect 9600 -910 10430 -810
rect 7650 -1140 7810 -990
rect 4890 -1300 5000 -1210
rect 5000 -1300 5120 -1210
rect 6890 -1300 7000 -1210
rect 7000 -1300 7120 -1210
rect 7935 -1285 8005 -1215
rect 8460 -1060 8550 -1050
rect 8460 -1210 8480 -1060
rect 8480 -1210 8530 -1060
rect 8530 -1210 8550 -1060
rect 2110 -1400 2220 -1340
rect 2620 -1400 2730 -1340
rect 2370 -1580 2550 -1550
rect 2880 -1580 3060 -1550
rect 9590 -1060 9680 -1050
rect 9590 -1210 9610 -1060
rect 9610 -1210 9660 -1060
rect 9660 -1210 9680 -1060
rect 8630 -1320 8710 -1240
rect 9760 -1320 9840 -1240
rect 3250 -1580 4810 -1550
rect 5250 -1580 5260 -1540
rect 5260 -1580 6800 -1540
rect 6800 -1580 6810 -1540
rect 2110 -1640 8480 -1580
rect 8480 -1640 8530 -1580
rect 8530 -1640 11010 -1580
rect 2110 -2150 11010 -1640
<< metal1 >>
rect 7150 -200 8150 -180
rect 860 -240 1930 -220
rect 860 -710 880 -240
rect 1910 -710 1930 -240
rect 7150 -370 7170 -200
rect 8130 -370 8150 -200
rect 7150 -380 8150 -370
rect 8350 -200 9350 -180
rect 8350 -370 8370 -200
rect 9330 -370 9350 -200
rect 8350 -380 9350 -370
rect 9480 -200 10480 -180
rect 9480 -370 9500 -200
rect 10460 -370 10480 -200
rect 9480 -380 10480 -370
rect 10620 -394 10850 -380
rect 10620 -400 10636 -394
rect 10620 -600 10630 -400
rect 10620 -606 10636 -600
rect 10836 -606 10850 -394
rect 10620 -620 10850 -606
rect 7250 -640 8120 -620
rect 860 -740 1090 -710
rect 1190 -740 1930 -710
rect 860 -750 1930 -740
rect 2360 -680 2560 -674
rect 820 -1050 1220 -1040
rect 820 -1120 840 -1050
rect 1200 -1120 1220 -1050
rect 820 -1130 1220 -1120
rect 1450 -1050 1930 -1040
rect 1450 -1120 1460 -1050
rect 1910 -1120 1930 -1050
rect 1450 -1130 1930 -1120
rect 2360 -1090 2560 -880
rect 2360 -1130 2380 -1090
rect 2540 -1130 2560 -1090
rect 2360 -1150 2560 -1130
rect 2870 -680 3070 -674
rect 2870 -1090 3070 -880
rect 3230 -800 4830 -790
rect 3230 -900 3250 -800
rect 4810 -900 4830 -800
rect 3230 -910 4830 -900
rect 5230 -800 6830 -790
rect 5230 -900 5250 -800
rect 6810 -900 6830 -800
rect 5230 -910 6830 -900
rect 7250 -910 7270 -640
rect 8100 -910 8120 -640
rect 7250 -920 8120 -910
rect 8450 -640 9320 -620
rect 8450 -910 8470 -640
rect 9300 -910 9320 -640
rect 8450 -920 9320 -910
rect 9580 -640 10450 -620
rect 9580 -910 9600 -640
rect 10430 -910 10450 -640
rect 9580 -920 10450 -910
rect 2870 -1140 2890 -1090
rect 3050 -1140 3070 -1090
rect 2870 -1150 3070 -1140
rect 7630 -990 7830 -920
rect 7630 -1140 7650 -990
rect 7810 -994 7830 -990
rect 7816 -1134 7830 -994
rect 7810 -1140 7830 -1134
rect 7630 -1200 7830 -1140
rect 8450 -1050 8560 -920
rect 4860 -1210 5150 -1200
rect 4860 -1300 4890 -1210
rect 5130 -1300 5150 -1210
rect 4860 -1310 5150 -1300
rect 6860 -1210 7150 -1200
rect 6860 -1300 6890 -1210
rect 7130 -1300 7150 -1210
rect 7923 -1215 8017 -1209
rect 7923 -1221 7935 -1215
rect 8005 -1221 8017 -1215
rect 7923 -1291 7929 -1221
rect 8011 -1291 8017 -1221
rect 8450 -1210 8460 -1050
rect 8550 -1210 8560 -1050
rect 8450 -1230 8560 -1210
rect 9580 -1050 9690 -920
rect 9580 -1210 9590 -1050
rect 9680 -1210 9690 -1050
rect 8618 -1240 8722 -1234
rect 9580 -1240 9690 -1210
rect 9748 -1240 9852 -1234
rect 8618 -1246 8630 -1240
rect 8710 -1246 8722 -1240
rect 7929 -1297 8011 -1291
rect 6860 -1310 7150 -1300
rect 8618 -1326 8624 -1246
rect 8716 -1326 8722 -1246
rect 9748 -1246 9760 -1240
rect 9840 -1246 9852 -1240
rect 9748 -1326 9754 -1246
rect 9846 -1326 9852 -1246
rect 2090 -1340 2310 -1330
rect 2090 -1400 2100 -1340
rect 2280 -1400 2310 -1340
rect 2090 -1410 2310 -1400
rect 2600 -1340 2820 -1330
rect 8624 -1332 8716 -1326
rect 9754 -1332 9846 -1326
rect 2600 -1400 2610 -1340
rect 2790 -1400 2820 -1340
rect 2600 -1410 2820 -1400
rect 1530 -1540 11030 -1530
rect 1530 -1550 5250 -1540
rect 1530 -1580 2370 -1550
rect 2550 -1580 2880 -1550
rect 3060 -1580 3250 -1550
rect 4810 -1580 5250 -1550
rect 6810 -1580 11030 -1540
rect 1530 -2150 2110 -1580
rect 11010 -2150 11030 -1580
rect 1530 -2170 11030 -2150
<< via1 >>
rect 880 -710 1910 -240
rect 7170 -370 8130 -200
rect 8370 -370 9330 -200
rect 9500 -370 10460 -200
rect 10636 -400 10836 -394
rect 10636 -600 10830 -400
rect 10830 -600 10836 -400
rect 10636 -606 10836 -600
rect 2360 -880 2560 -680
rect 840 -1120 1110 -1050
rect 1110 -1120 1200 -1050
rect 1460 -1120 1470 -1050
rect 1470 -1120 1580 -1050
rect 1580 -1120 1910 -1050
rect 2870 -880 3070 -680
rect 3250 -810 4810 -800
rect 3250 -900 4810 -810
rect 5250 -810 6810 -800
rect 5250 -900 6810 -810
rect 7270 -910 8100 -640
rect 8470 -910 9300 -640
rect 9600 -910 10430 -640
rect 7650 -1140 7810 -990
rect 7810 -1134 7816 -994
rect 4890 -1300 5120 -1210
rect 5120 -1300 5130 -1210
rect 6890 -1300 7120 -1210
rect 7120 -1300 7130 -1210
rect 7929 -1285 7935 -1221
rect 7935 -1285 8005 -1221
rect 8005 -1285 8011 -1221
rect 7929 -1291 8011 -1285
rect 8460 -1210 8550 -1050
rect 9590 -1210 9680 -1050
rect 8624 -1320 8630 -1246
rect 8630 -1320 8710 -1246
rect 8710 -1320 8716 -1246
rect 8624 -1326 8716 -1320
rect 9754 -1320 9760 -1246
rect 9760 -1320 9840 -1246
rect 9840 -1320 9846 -1246
rect 9754 -1326 9846 -1320
rect 2100 -1400 2110 -1340
rect 2110 -1400 2220 -1340
rect 2220 -1400 2280 -1340
rect 2610 -1400 2620 -1340
rect 2620 -1400 2730 -1340
rect 2730 -1400 2790 -1340
<< metal2 >>
rect 7150 -200 8150 -180
rect 860 -240 1930 -220
rect 860 -710 880 -240
rect 1910 -710 1930 -240
rect 7150 -370 7170 -200
rect 8130 -370 8150 -200
rect 7150 -380 8150 -370
rect 8350 -200 9350 -180
rect 8350 -370 8370 -200
rect 9330 -370 9350 -200
rect 8350 -380 9350 -370
rect 9480 -200 10480 -180
rect 9480 -370 9500 -200
rect 10460 -370 10480 -200
rect 9480 -380 10480 -370
rect 10620 -394 10850 -380
rect 10620 -606 10636 -394
rect 10836 -606 10850 -394
rect 10620 -620 10850 -606
rect 7250 -640 8120 -620
rect 860 -750 1930 -710
rect 2350 -680 2570 -670
rect 2350 -880 2360 -680
rect 2560 -880 2570 -680
rect 2350 -890 2570 -880
rect 2860 -680 3080 -670
rect 2860 -880 2870 -680
rect 3070 -880 3080 -680
rect 2860 -890 3080 -880
rect 3230 -800 4830 -790
rect 3230 -900 3250 -800
rect 4810 -900 4830 -800
rect 3230 -910 4830 -900
rect 5230 -800 6830 -790
rect 5230 -900 5250 -800
rect 6810 -900 6830 -800
rect 5230 -910 6830 -900
rect 7250 -910 7270 -640
rect 8100 -910 8120 -640
rect 7250 -920 8120 -910
rect 8450 -640 9320 -620
rect 8450 -910 8470 -640
rect 9300 -910 9320 -640
rect 8450 -920 9320 -910
rect 9580 -640 10450 -620
rect 9580 -910 9600 -640
rect 10430 -910 10450 -640
rect 9580 -920 10450 -910
rect 7630 -990 7830 -920
rect 790 -1050 1220 -1040
rect 790 -1120 840 -1050
rect 1200 -1120 1220 -1050
rect 790 -1130 1220 -1120
rect 1450 -1050 1930 -1040
rect 1450 -1120 1460 -1050
rect 1910 -1120 1930 -1050
rect 1450 -1130 1930 -1120
rect 7630 -1140 7650 -990
rect 7810 -994 7830 -990
rect 7816 -1134 7830 -994
rect 7810 -1140 7830 -1134
rect 7630 -1200 7830 -1140
rect 8450 -1050 8560 -920
rect 4860 -1210 5150 -1200
rect 4860 -1300 4890 -1210
rect 5130 -1300 5150 -1210
rect 4860 -1310 5150 -1300
rect 6860 -1210 7150 -1200
rect 8450 -1210 8460 -1050
rect 8550 -1210 8560 -1050
rect 6860 -1300 6890 -1210
rect 7130 -1300 7150 -1210
rect 7930 -1221 8010 -1210
rect 7923 -1291 7929 -1221
rect 8011 -1291 8017 -1221
rect 8450 -1230 8560 -1210
rect 9580 -1050 9690 -920
rect 9580 -1210 9590 -1050
rect 9680 -1210 9690 -1050
rect 9580 -1240 9690 -1210
rect 6860 -1310 7150 -1300
rect 2090 -1340 2310 -1330
rect 2090 -1400 2100 -1340
rect 2280 -1400 2310 -1340
rect 2090 -1410 2310 -1400
rect 2600 -1340 2820 -1330
rect 2600 -1400 2610 -1340
rect 2790 -1400 2820 -1340
rect 2600 -1410 2820 -1400
rect 2090 -2235 2180 -1410
rect 2600 -2225 2690 -1410
rect 5040 -2205 5150 -1310
rect 7040 -2205 7150 -1310
rect 7930 -2230 8010 -1291
rect 8618 -1326 8624 -1246
rect 8716 -1326 8722 -1246
rect 9748 -1326 9754 -1246
rect 9846 -1326 9852 -1246
rect 8630 -2240 8710 -1326
rect 9760 -2240 9840 -1326
<< via2 >>
rect 7170 -370 8130 -200
rect 8370 -370 9330 -200
rect 9500 -370 10460 -200
rect 10636 -606 10836 -394
rect 2360 -880 2560 -680
rect 2870 -880 3070 -680
rect 3250 -900 4810 -800
rect 5250 -900 6810 -800
rect 7270 -910 8100 -640
rect 8470 -910 9300 -640
rect 9600 -910 10430 -640
rect 1470 -1120 1910 -1050
rect 7664 -1134 7816 -1040
rect 8460 -1210 8550 -1050
rect 9590 -1210 9680 -1050
<< metal3 >>
rect 7150 -200 8150 -60
rect 7150 -370 7170 -200
rect 8130 -370 8150 -200
rect 2360 -670 2560 -370
rect 2870 -670 3070 -370
rect 7150 -380 8150 -370
rect 8350 -200 9350 -60
rect 8350 -370 8370 -200
rect 9330 -370 9350 -200
rect 8350 -380 9350 -370
rect 9480 -200 10480 -60
rect 9480 -370 9500 -200
rect 10460 -370 10480 -200
rect 9480 -380 10480 -370
rect 10620 -394 10850 -380
rect 10620 -606 10636 -394
rect 10836 -400 10850 -394
rect 10836 -600 11230 -400
rect 10836 -606 10850 -600
rect 10620 -620 10850 -606
rect 7250 -640 8120 -620
rect 2350 -680 2570 -670
rect 2350 -880 2360 -680
rect 2560 -880 2570 -680
rect 2350 -890 2570 -880
rect 2860 -680 3080 -670
rect 2860 -880 2870 -680
rect 3070 -880 3080 -680
rect 2860 -890 3080 -880
rect 3230 -800 4830 -680
rect 3230 -900 3250 -800
rect 4810 -900 4830 -800
rect 3230 -910 4830 -900
rect 5230 -800 6830 -680
rect 5230 -900 5250 -800
rect 6810 -900 6830 -800
rect 5230 -910 6830 -900
rect 7250 -910 7270 -640
rect 8100 -910 8120 -640
rect 7250 -920 8120 -910
rect 8450 -640 9320 -620
rect 8450 -910 8470 -640
rect 9300 -910 9320 -640
rect 8450 -920 9320 -910
rect 9580 -640 10450 -620
rect 9580 -910 9600 -640
rect 10430 -910 10450 -640
rect 9580 -920 10450 -910
rect 7630 -1040 7830 -920
rect 1450 -1050 1930 -1040
rect 1450 -1120 1470 -1050
rect 1910 -1120 1930 -1050
rect 1450 -1130 1930 -1120
rect 1840 -2236 1930 -1130
rect 7630 -1134 7664 -1040
rect 7816 -1134 7830 -1040
rect 7630 -1150 7830 -1134
rect 8450 -1050 8560 -920
rect 8450 -1210 8460 -1050
rect 8550 -1210 8560 -1050
rect 8450 -1230 8560 -1210
rect 9580 -1050 9690 -920
rect 9580 -1210 9590 -1050
rect 9680 -1210 9690 -1050
rect 9580 -1230 9690 -1210
<< labels >>
rlabel metal1 870 -670 870 -670 1 VDD
port 1 n
rlabel metal2 2130 -1630 2130 -1630 1 NB1
port 4 n
rlabel metal2 2640 -1630 2640 -1630 1 NB2
port 5 n
rlabel metal2 5090 -1630 5090 -1630 1 OUT_IB
port 6 n
rlabel metal2 7100 -1630 7100 -1630 1 AMP_IB
port 7 n
rlabel metal1 1650 -1540 1650 -1540 1 GND
port 12 n
rlabel metal3 1840 -2236 1930 -2200 1 SF_IB
port 13 n
rlabel metal2 8670 -2200 8670 -2200 1 BIAS1_OUT
port 14 n
rlabel metal2 7970 -2190 7970 -2190 1 BIAS2_OUT
port 15 n
rlabel metal3 8680 -90 8680 -90 1 BIAS1
port 17 n
rlabel metal3 7480 -100 7480 -100 1 BIAS2
port 18 n
rlabel metal3 11220 -500 11220 -500 1 ADC_ON
port 16 n
rlabel metal2 9800 -2200 9800 -2200 1 SA_IREF_OUT
port 19 n
rlabel metal3 9800 -90 9800 -90 1 SA_IREF
port 20 n
<< end >>
