magic
tech sky130B
magscale 1 2
timestamp 1608351071
<< pwell >>
rect -211 -208 211 208
<< nmos >>
rect -15 -60 15 60
<< ndiff >>
rect -73 48 -15 60
rect -73 -48 -61 48
rect -27 -48 -15 48
rect -73 -60 -15 -48
rect 15 48 73 60
rect 15 -48 27 48
rect 61 -48 73 48
rect 15 -60 73 -48
<< ndiffc >>
rect -61 -48 -27 48
rect 27 -48 61 48
<< psubdiff >>
rect -175 76 -141 138
rect 141 76 175 138
rect -175 -138 -141 -76
rect 141 -138 175 -76
rect -175 -172 -79 -138
rect 79 -172 175 -138
<< psubdiffcont >>
rect -175 -76 -141 76
rect 141 -76 175 76
rect -79 -172 79 -138
<< poly >>
rect -15 60 15 86
rect -15 -86 15 -60
<< locali >>
rect -175 138 175 172
rect -175 76 -141 138
rect 141 76 175 138
rect -61 48 -27 64
rect -61 -64 -27 -48
rect 27 48 61 64
rect 27 -64 61 -48
rect -175 -138 -141 -76
rect 141 -138 175 -76
rect -175 -172 -79 -138
rect 79 -172 175 -138
<< viali >>
rect -61 -48 -27 48
rect 27 -48 61 48
<< metal1 >>
rect -67 48 -21 60
rect -67 -48 -61 48
rect -27 -48 -21 48
rect -67 -60 -21 -48
rect 21 48 67 60
rect 21 -48 27 48
rect 61 -48 67 48
rect 21 -60 67 -48
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -158 -155 158 155
string parameters w 0.6 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
