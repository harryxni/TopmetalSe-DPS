magic
tech sky130B
magscale 1 2
timestamp 1608325973
<< nwell >>
rect -97 -60 503 767
<< pwell >>
rect -112 -910 511 -158
<< psubdiff >>
rect -51 -679 461 -615
rect -51 -850 -25 -679
rect 434 -850 461 -679
rect -51 -851 461 -850
<< nsubdiff >>
rect -45 502 459 726
<< psubdiffcont >>
rect -25 -850 434 -679
<< locali >>
rect -33 725 451 726
rect -41 -850 -25 -849
rect 434 -850 450 -849
<< viali >>
rect -48 500 459 725
rect -54 -679 461 -618
rect -54 -849 -25 -679
rect -25 -849 434 -679
rect 434 -849 461 -679
<< metal1 >>
rect -60 725 471 731
rect -60 500 -48 725
rect 459 500 471 725
rect -60 494 471 500
rect -128 297 -118 443
rect -36 438 -26 443
rect -36 383 289 438
rect -36 297 -26 383
rect 63 165 73 347
rect 128 165 138 347
rect 174 166 184 347
rect 236 166 246 347
rect 278 164 288 346
rect 343 164 353 346
rect -233 21 -223 164
rect -143 127 -133 164
rect -143 72 226 127
rect -143 21 -133 72
rect -119 -349 -109 -209
rect -50 -290 -40 -209
rect -50 -345 282 -290
rect -50 -349 -40 -345
rect -267 -447 127 -392
rect 264 -489 274 -382
rect 341 -489 351 -382
rect -238 -638 -228 -495
rect -124 -550 184 -495
rect -124 -638 -114 -550
rect -66 -618 473 -612
rect -66 -849 -54 -618
rect 461 -849 473 -618
rect -66 -855 473 -849
<< via1 >>
rect -48 500 459 725
rect -118 297 -36 443
rect 73 165 128 347
rect 184 166 236 347
rect 288 164 343 346
rect -223 21 -143 164
rect -109 -349 -50 -209
rect 274 -489 341 -382
rect -228 -638 -124 -495
<< metal2 >>
rect -48 725 459 735
rect -48 490 459 500
rect -118 443 -36 453
rect 74 357 125 358
rect 182 357 235 490
rect -118 287 -36 297
rect 73 347 128 357
rect -223 164 -143 174
rect -223 11 -143 21
rect -211 -485 -155 11
rect -110 -199 -54 287
rect 73 155 128 165
rect 182 347 236 357
rect 182 166 184 347
rect 182 156 236 166
rect 288 346 343 356
rect 74 82 125 155
rect 288 154 343 164
rect 291 82 342 154
rect 74 31 342 82
rect -110 -209 -50 -199
rect -110 -349 -109 -209
rect -110 -350 -50 -349
rect -109 -359 -50 -350
rect 291 -372 342 31
rect 274 -382 342 -372
rect -228 -495 -124 -485
rect 341 -489 342 -382
rect 274 -496 342 -489
rect 274 -499 341 -496
rect -228 -648 -124 -638
use sky130_fd_pr__pfet_01v8_H49BFK  sky130_fd_pr__pfet_01v8_H49BFK_0
timestamp 1608325295
transform 1 0 210 0 1 256
box -263 -309 263 309
use sky130_fd_pr__nfet_01v8_TFZGL8  sky130_fd_pr__nfet_01v8_TFZGL8_0
timestamp 1608325973
transform 1 0 201 0 1 -421
box -263 -255 263 255
<< labels >>
rlabel metal1 -98 383 289 438 1 A
rlabel nwell -48 500 459 725 1 vdd
rlabel metal1 -233 21 -223 164 1 B
rlabel metal1 -128 297 -118 443 1 A
rlabel pwell -54 -849 461 -618 1 bulk_n
rlabel space -267 -447 128 -392 1 vss
rlabel metal2 291 -382 342 164 1 out
<< end >>
