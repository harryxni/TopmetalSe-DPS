magic
tech sky130B
magscale 1 2
timestamp 1662181890
<< metal1 >>
rect -1895 3270 -1745 3276
rect -600 3270 -210 3320
rect -1745 3120 420 3270
rect -1895 3114 -1745 3120
rect -600 2890 -210 3120
rect -81 330 -75 480
rect 75 330 420 480
<< via1 >>
rect -1895 3120 -1745 3270
rect -75 330 75 480
<< metal2 >>
rect -2820 3048 -2680 3450
rect -2820 2992 -2778 3048
rect -2722 2992 -2680 3048
rect -2820 -70 -2680 2992
rect -2310 2848 -2170 3490
rect -1895 3270 -1745 3279
rect -1901 3120 -1895 3270
rect -1745 3120 -1739 3270
rect -1895 3111 -1745 3120
rect -2310 2792 -2268 2848
rect -2212 2792 -2170 2848
rect -2310 -90 -2170 2792
rect -1431 2548 -1328 2610
rect -1431 2492 -1408 2548
rect -1352 2492 -1328 2548
rect -1431 1970 -1328 2492
rect -920 738 -780 870
rect -920 682 -878 738
rect -822 682 -780 738
rect -920 500 -780 682
rect -75 480 75 486
rect -84 330 -75 480
rect 75 330 84 480
rect -75 324 75 330
<< via2 >>
rect -2778 2992 -2722 3048
rect -1895 3120 -1745 3270
rect -2268 2792 -2212 2848
rect -1408 2492 -1352 2548
rect -878 682 -822 738
rect -75 330 75 480
<< metal3 >>
rect -1900 3275 -1740 3281
rect -1900 3120 -1895 3125
rect -1745 3120 -1740 3125
rect -1900 3115 -1740 3120
rect -2783 3050 -2717 3053
rect -2783 3048 250 3050
rect -2783 2992 -2778 3048
rect -2722 2992 250 3048
rect -2783 2990 250 2992
rect -2783 2987 -2717 2990
rect -2273 2850 -2207 2853
rect -2273 2848 60 2850
rect -2273 2792 -2268 2848
rect -2212 2792 60 2848
rect -2273 2790 60 2792
rect -2273 2787 -2207 2790
rect -1413 2550 -1347 2553
rect -1413 2548 160 2550
rect -1413 2492 -1408 2548
rect -1352 2492 160 2548
rect -1413 2490 160 2492
rect -1413 2487 -1347 2490
rect -883 740 -817 743
rect -883 738 80 740
rect -883 682 -878 738
rect -822 682 80 738
rect -883 680 80 682
rect -883 677 -817 680
rect -475 480 -325 486
rect -80 480 80 485
rect -325 330 -75 480
rect 75 330 80 480
rect -475 324 -325 330
rect -80 325 80 330
<< via3 >>
rect -1900 3270 -1740 3275
rect -1900 3125 -1895 3270
rect -1895 3125 -1745 3270
rect -1745 3125 -1740 3270
rect -475 330 -325 480
<< metal4 >>
rect -2010 3275 -1620 3630
rect -2010 3125 -1900 3275
rect -1740 3125 -1620 3275
rect -610 3160 -220 3640
rect -2010 3120 -1620 3125
rect -580 3030 -230 3160
<< via4 >>
rect -1980 170 -1650 3060
rect -560 480 -240 3030
rect -560 330 -475 480
rect -475 330 -325 480
rect -325 330 -240 480
rect -560 170 -240 330
<< metal5 >>
rect -2010 3060 -1620 3630
rect -2010 170 -1980 3060
rect -1650 170 -1620 3060
rect -2010 -130 -1620 170
rect -610 3320 -220 3640
rect -610 3030 -210 3320
rect -610 170 -560 3030
rect -240 170 -210 3030
rect -610 -120 -210 170
use pixel  pixel_0
timestamp 1662180122
transform 1 0 470 0 1 3000
box -470 -3000 3090 570
<< end >>
