** sch_path: /home/hni/topmetal_dps/xschem/sens_amp.sch
**.subckt sens_amp REF V_IN OUT SA_IREF
*.ipin REF
*.ipin V_IN
*.opin OUT
*.ipin SA_IREF
XM5 net1 GN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1
XM6 GN GN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1
XM23 net1 V_IN net2 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1
XM16 GN REF net2 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1
XM1 OUT net1 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=3 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 SA_IREF GND GND sky130_fd_pr__nfet_01v8_lvt L=1 W=0.5 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1
**.ends
.GLOBAL GND
.end
