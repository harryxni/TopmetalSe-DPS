magic
tech sky130B
magscale 1 2
timestamp 1608322001
<< error_p >>
rect -29 181 29 187
rect -29 147 -17 181
rect -29 141 29 147
<< pwell >>
rect -211 -319 211 319
<< nmos >>
rect -15 -109 15 109
<< ndiff >>
rect -73 97 -15 109
rect -73 -97 -61 97
rect -27 -97 -15 97
rect -73 -109 -15 -97
rect 15 97 73 109
rect 15 -97 27 97
rect 61 -97 73 97
rect 15 -109 73 -97
<< ndiffc >>
rect -61 -97 -27 97
rect 27 -97 61 97
<< psubdiff >>
rect -175 249 -79 283
rect 79 249 175 283
rect -175 187 -141 249
rect 141 187 175 249
rect -175 -249 -141 -187
rect 141 -249 175 -187
rect -175 -283 -79 -249
rect 79 -283 175 -249
<< psubdiffcont >>
rect -79 249 79 283
rect -175 -187 -141 187
rect 141 -187 175 187
rect -79 -283 79 -249
<< poly >>
rect -33 181 33 197
rect -33 147 -17 181
rect 17 147 33 181
rect -33 131 33 147
rect -15 109 15 131
rect -15 -143 15 -109
<< polycont >>
rect -17 147 17 181
<< locali >>
rect -175 249 -79 283
rect 79 249 175 283
rect -175 187 -141 249
rect 141 187 175 249
rect -33 147 -17 181
rect 17 147 33 181
rect -61 97 -27 113
rect -61 -113 -27 -97
rect 27 97 61 113
rect 27 -113 61 -97
rect -175 -249 -141 -187
rect 141 -249 175 -187
rect -175 -283 -79 -249
rect 79 -283 175 -249
<< viali >>
rect -17 147 17 181
rect -61 -97 -27 97
rect 27 -97 61 97
<< metal1 >>
rect -29 181 29 187
rect -29 147 -17 181
rect 17 147 29 181
rect -29 141 29 147
rect -67 97 -21 109
rect -67 -97 -61 97
rect -27 -97 -21 97
rect -67 -109 -21 -97
rect 21 97 67 109
rect 21 -97 27 97
rect 61 -97 67 97
rect 21 -109 67 -97
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -158 -266 158 266
string parameters w 1.09 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
