magic
tech sky130B
magscale 1 2
timestamp 1606423877
<< error_p >>
rect -560 1217 -502 1223
rect -442 1217 -384 1223
rect -324 1217 -266 1223
rect -206 1217 -148 1223
rect -88 1217 -30 1223
rect 30 1217 88 1223
rect 148 1217 206 1223
rect 266 1217 324 1223
rect 384 1217 442 1223
rect 502 1217 560 1223
rect -560 1183 -548 1217
rect -442 1183 -430 1217
rect -324 1183 -312 1217
rect -206 1183 -194 1217
rect -88 1183 -76 1217
rect 30 1183 42 1217
rect 148 1183 160 1217
rect 266 1183 278 1217
rect 384 1183 396 1217
rect 502 1183 514 1217
rect -560 1177 -502 1183
rect -442 1177 -384 1183
rect -324 1177 -266 1183
rect -206 1177 -148 1183
rect -88 1177 -30 1183
rect 30 1177 88 1183
rect 148 1177 206 1183
rect 266 1177 324 1183
rect 384 1177 442 1183
rect 502 1177 560 1183
rect -560 489 -502 495
rect -442 489 -384 495
rect -324 489 -266 495
rect -206 489 -148 495
rect -88 489 -30 495
rect 30 489 88 495
rect 148 489 206 495
rect 266 489 324 495
rect 384 489 442 495
rect 502 489 560 495
rect -560 455 -548 489
rect -442 455 -430 489
rect -324 455 -312 489
rect -206 455 -194 489
rect -88 455 -76 489
rect 30 455 42 489
rect 148 455 160 489
rect 266 455 278 489
rect 384 455 396 489
rect 502 455 514 489
rect -560 449 -502 455
rect -442 449 -384 455
rect -324 449 -266 455
rect -206 449 -148 455
rect -88 449 -30 455
rect 30 449 88 455
rect 148 449 206 455
rect 266 449 324 455
rect 384 449 442 455
rect 502 449 560 455
rect -560 381 -502 387
rect -442 381 -384 387
rect -324 381 -266 387
rect -206 381 -148 387
rect -88 381 -30 387
rect 30 381 88 387
rect 148 381 206 387
rect 266 381 324 387
rect 384 381 442 387
rect 502 381 560 387
rect -560 347 -548 381
rect -442 347 -430 381
rect -324 347 -312 381
rect -206 347 -194 381
rect -88 347 -76 381
rect 30 347 42 381
rect 148 347 160 381
rect 266 347 278 381
rect 384 347 396 381
rect 502 347 514 381
rect -560 341 -502 347
rect -442 341 -384 347
rect -324 341 -266 347
rect -206 341 -148 347
rect -88 341 -30 347
rect 30 341 88 347
rect 148 341 206 347
rect 266 341 324 347
rect 384 341 442 347
rect 502 341 560 347
rect -560 -347 -502 -341
rect -442 -347 -384 -341
rect -324 -347 -266 -341
rect -206 -347 -148 -341
rect -88 -347 -30 -341
rect 30 -347 88 -341
rect 148 -347 206 -341
rect 266 -347 324 -341
rect 384 -347 442 -341
rect 502 -347 560 -341
rect -560 -381 -548 -347
rect -442 -381 -430 -347
rect -324 -381 -312 -347
rect -206 -381 -194 -347
rect -88 -381 -76 -347
rect 30 -381 42 -347
rect 148 -381 160 -347
rect 266 -381 278 -347
rect 384 -381 396 -347
rect 502 -381 514 -347
rect -560 -387 -502 -381
rect -442 -387 -384 -381
rect -324 -387 -266 -381
rect -206 -387 -148 -381
rect -88 -387 -30 -381
rect 30 -387 88 -381
rect 148 -387 206 -381
rect 266 -387 324 -381
rect 384 -387 442 -381
rect 502 -387 560 -381
rect -560 -455 -502 -449
rect -442 -455 -384 -449
rect -324 -455 -266 -449
rect -206 -455 -148 -449
rect -88 -455 -30 -449
rect 30 -455 88 -449
rect 148 -455 206 -449
rect 266 -455 324 -449
rect 384 -455 442 -449
rect 502 -455 560 -449
rect -560 -489 -548 -455
rect -442 -489 -430 -455
rect -324 -489 -312 -455
rect -206 -489 -194 -455
rect -88 -489 -76 -455
rect 30 -489 42 -455
rect 148 -489 160 -455
rect 266 -489 278 -455
rect 384 -489 396 -455
rect 502 -489 514 -455
rect -560 -495 -502 -489
rect -442 -495 -384 -489
rect -324 -495 -266 -489
rect -206 -495 -148 -489
rect -88 -495 -30 -489
rect 30 -495 88 -489
rect 148 -495 206 -489
rect 266 -495 324 -489
rect 384 -495 442 -489
rect 502 -495 560 -489
rect -560 -1183 -502 -1177
rect -442 -1183 -384 -1177
rect -324 -1183 -266 -1177
rect -206 -1183 -148 -1177
rect -88 -1183 -30 -1177
rect 30 -1183 88 -1177
rect 148 -1183 206 -1177
rect 266 -1183 324 -1177
rect 384 -1183 442 -1177
rect 502 -1183 560 -1177
rect -560 -1217 -548 -1183
rect -442 -1217 -430 -1183
rect -324 -1217 -312 -1183
rect -206 -1217 -194 -1183
rect -88 -1217 -76 -1183
rect 30 -1217 42 -1183
rect 148 -1217 160 -1183
rect 266 -1217 278 -1183
rect 384 -1217 396 -1183
rect 502 -1217 514 -1183
rect -560 -1223 -502 -1217
rect -442 -1223 -384 -1217
rect -324 -1223 -266 -1217
rect -206 -1223 -148 -1217
rect -88 -1223 -30 -1217
rect 30 -1223 88 -1217
rect 148 -1223 206 -1217
rect 266 -1223 324 -1217
rect 384 -1223 442 -1217
rect 502 -1223 560 -1217
<< nwell >>
rect -757 -1355 757 1355
<< pmos >>
rect -561 536 -501 1136
rect -443 536 -383 1136
rect -325 536 -265 1136
rect -207 536 -147 1136
rect -89 536 -29 1136
rect 29 536 89 1136
rect 147 536 207 1136
rect 265 536 325 1136
rect 383 536 443 1136
rect 501 536 561 1136
rect -561 -300 -501 300
rect -443 -300 -383 300
rect -325 -300 -265 300
rect -207 -300 -147 300
rect -89 -300 -29 300
rect 29 -300 89 300
rect 147 -300 207 300
rect 265 -300 325 300
rect 383 -300 443 300
rect 501 -300 561 300
rect -561 -1136 -501 -536
rect -443 -1136 -383 -536
rect -325 -1136 -265 -536
rect -207 -1136 -147 -536
rect -89 -1136 -29 -536
rect 29 -1136 89 -536
rect 147 -1136 207 -536
rect 265 -1136 325 -536
rect 383 -1136 443 -536
rect 501 -1136 561 -536
<< pdiff >>
rect -619 1124 -561 1136
rect -619 548 -607 1124
rect -573 548 -561 1124
rect -619 536 -561 548
rect -501 1124 -443 1136
rect -501 548 -489 1124
rect -455 548 -443 1124
rect -501 536 -443 548
rect -383 1124 -325 1136
rect -383 548 -371 1124
rect -337 548 -325 1124
rect -383 536 -325 548
rect -265 1124 -207 1136
rect -265 548 -253 1124
rect -219 548 -207 1124
rect -265 536 -207 548
rect -147 1124 -89 1136
rect -147 548 -135 1124
rect -101 548 -89 1124
rect -147 536 -89 548
rect -29 1124 29 1136
rect -29 548 -17 1124
rect 17 548 29 1124
rect -29 536 29 548
rect 89 1124 147 1136
rect 89 548 101 1124
rect 135 548 147 1124
rect 89 536 147 548
rect 207 1124 265 1136
rect 207 548 219 1124
rect 253 548 265 1124
rect 207 536 265 548
rect 325 1124 383 1136
rect 325 548 337 1124
rect 371 548 383 1124
rect 325 536 383 548
rect 443 1124 501 1136
rect 443 548 455 1124
rect 489 548 501 1124
rect 443 536 501 548
rect 561 1124 619 1136
rect 561 548 573 1124
rect 607 548 619 1124
rect 561 536 619 548
rect -619 288 -561 300
rect -619 -288 -607 288
rect -573 -288 -561 288
rect -619 -300 -561 -288
rect -501 288 -443 300
rect -501 -288 -489 288
rect -455 -288 -443 288
rect -501 -300 -443 -288
rect -383 288 -325 300
rect -383 -288 -371 288
rect -337 -288 -325 288
rect -383 -300 -325 -288
rect -265 288 -207 300
rect -265 -288 -253 288
rect -219 -288 -207 288
rect -265 -300 -207 -288
rect -147 288 -89 300
rect -147 -288 -135 288
rect -101 -288 -89 288
rect -147 -300 -89 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 89 288 147 300
rect 89 -288 101 288
rect 135 -288 147 288
rect 89 -300 147 -288
rect 207 288 265 300
rect 207 -288 219 288
rect 253 -288 265 288
rect 207 -300 265 -288
rect 325 288 383 300
rect 325 -288 337 288
rect 371 -288 383 288
rect 325 -300 383 -288
rect 443 288 501 300
rect 443 -288 455 288
rect 489 -288 501 288
rect 443 -300 501 -288
rect 561 288 619 300
rect 561 -288 573 288
rect 607 -288 619 288
rect 561 -300 619 -288
rect -619 -548 -561 -536
rect -619 -1124 -607 -548
rect -573 -1124 -561 -548
rect -619 -1136 -561 -1124
rect -501 -548 -443 -536
rect -501 -1124 -489 -548
rect -455 -1124 -443 -548
rect -501 -1136 -443 -1124
rect -383 -548 -325 -536
rect -383 -1124 -371 -548
rect -337 -1124 -325 -548
rect -383 -1136 -325 -1124
rect -265 -548 -207 -536
rect -265 -1124 -253 -548
rect -219 -1124 -207 -548
rect -265 -1136 -207 -1124
rect -147 -548 -89 -536
rect -147 -1124 -135 -548
rect -101 -1124 -89 -548
rect -147 -1136 -89 -1124
rect -29 -548 29 -536
rect -29 -1124 -17 -548
rect 17 -1124 29 -548
rect -29 -1136 29 -1124
rect 89 -548 147 -536
rect 89 -1124 101 -548
rect 135 -1124 147 -548
rect 89 -1136 147 -1124
rect 207 -548 265 -536
rect 207 -1124 219 -548
rect 253 -1124 265 -548
rect 207 -1136 265 -1124
rect 325 -548 383 -536
rect 325 -1124 337 -548
rect 371 -1124 383 -548
rect 325 -1136 383 -1124
rect 443 -548 501 -536
rect 443 -1124 455 -548
rect 489 -1124 501 -548
rect 443 -1136 501 -1124
rect 561 -548 619 -536
rect 561 -1124 573 -548
rect 607 -1124 619 -548
rect 561 -1136 619 -1124
<< pdiffc >>
rect -607 548 -573 1124
rect -489 548 -455 1124
rect -371 548 -337 1124
rect -253 548 -219 1124
rect -135 548 -101 1124
rect -17 548 17 1124
rect 101 548 135 1124
rect 219 548 253 1124
rect 337 548 371 1124
rect 455 548 489 1124
rect 573 548 607 1124
rect -607 -288 -573 288
rect -489 -288 -455 288
rect -371 -288 -337 288
rect -253 -288 -219 288
rect -135 -288 -101 288
rect -17 -288 17 288
rect 101 -288 135 288
rect 219 -288 253 288
rect 337 -288 371 288
rect 455 -288 489 288
rect 573 -288 607 288
rect -607 -1124 -573 -548
rect -489 -1124 -455 -548
rect -371 -1124 -337 -548
rect -253 -1124 -219 -548
rect -135 -1124 -101 -548
rect -17 -1124 17 -548
rect 101 -1124 135 -548
rect 219 -1124 253 -548
rect 337 -1124 371 -548
rect 455 -1124 489 -548
rect 573 -1124 607 -548
<< nsubdiff >>
rect -721 1285 -625 1319
rect 625 1285 721 1319
rect -721 1223 -687 1285
rect 687 1223 721 1285
rect -721 -1285 -687 -1223
rect 687 -1285 721 -1223
rect -721 -1319 -625 -1285
rect 625 -1319 721 -1285
<< nsubdiffcont >>
rect -625 1285 625 1319
rect -721 -1223 -687 1223
rect 687 -1223 721 1223
rect -625 -1319 625 -1285
<< poly >>
rect -564 1217 -498 1233
rect -564 1183 -548 1217
rect -514 1183 -498 1217
rect -564 1167 -498 1183
rect -446 1217 -380 1233
rect -446 1183 -430 1217
rect -396 1183 -380 1217
rect -446 1167 -380 1183
rect -328 1217 -262 1233
rect -328 1183 -312 1217
rect -278 1183 -262 1217
rect -328 1167 -262 1183
rect -210 1217 -144 1233
rect -210 1183 -194 1217
rect -160 1183 -144 1217
rect -210 1167 -144 1183
rect -92 1217 -26 1233
rect -92 1183 -76 1217
rect -42 1183 -26 1217
rect -92 1167 -26 1183
rect 26 1217 92 1233
rect 26 1183 42 1217
rect 76 1183 92 1217
rect 26 1167 92 1183
rect 144 1217 210 1233
rect 144 1183 160 1217
rect 194 1183 210 1217
rect 144 1167 210 1183
rect 262 1217 328 1233
rect 262 1183 278 1217
rect 312 1183 328 1217
rect 262 1167 328 1183
rect 380 1217 446 1233
rect 380 1183 396 1217
rect 430 1183 446 1217
rect 380 1167 446 1183
rect 498 1217 564 1233
rect 498 1183 514 1217
rect 548 1183 564 1217
rect 498 1167 564 1183
rect -561 1136 -501 1167
rect -443 1136 -383 1167
rect -325 1136 -265 1167
rect -207 1136 -147 1167
rect -89 1136 -29 1167
rect 29 1136 89 1167
rect 147 1136 207 1167
rect 265 1136 325 1167
rect 383 1136 443 1167
rect 501 1136 561 1167
rect -561 505 -501 536
rect -443 505 -383 536
rect -325 505 -265 536
rect -207 505 -147 536
rect -89 505 -29 536
rect 29 505 89 536
rect 147 505 207 536
rect 265 505 325 536
rect 383 505 443 536
rect 501 505 561 536
rect -564 489 -498 505
rect -564 455 -548 489
rect -514 455 -498 489
rect -564 439 -498 455
rect -446 489 -380 505
rect -446 455 -430 489
rect -396 455 -380 489
rect -446 439 -380 455
rect -328 489 -262 505
rect -328 455 -312 489
rect -278 455 -262 489
rect -328 439 -262 455
rect -210 489 -144 505
rect -210 455 -194 489
rect -160 455 -144 489
rect -210 439 -144 455
rect -92 489 -26 505
rect -92 455 -76 489
rect -42 455 -26 489
rect -92 439 -26 455
rect 26 489 92 505
rect 26 455 42 489
rect 76 455 92 489
rect 26 439 92 455
rect 144 489 210 505
rect 144 455 160 489
rect 194 455 210 489
rect 144 439 210 455
rect 262 489 328 505
rect 262 455 278 489
rect 312 455 328 489
rect 262 439 328 455
rect 380 489 446 505
rect 380 455 396 489
rect 430 455 446 489
rect 380 439 446 455
rect 498 489 564 505
rect 498 455 514 489
rect 548 455 564 489
rect 498 439 564 455
rect -564 381 -498 397
rect -564 347 -548 381
rect -514 347 -498 381
rect -564 331 -498 347
rect -446 381 -380 397
rect -446 347 -430 381
rect -396 347 -380 381
rect -446 331 -380 347
rect -328 381 -262 397
rect -328 347 -312 381
rect -278 347 -262 381
rect -328 331 -262 347
rect -210 381 -144 397
rect -210 347 -194 381
rect -160 347 -144 381
rect -210 331 -144 347
rect -92 381 -26 397
rect -92 347 -76 381
rect -42 347 -26 381
rect -92 331 -26 347
rect 26 381 92 397
rect 26 347 42 381
rect 76 347 92 381
rect 26 331 92 347
rect 144 381 210 397
rect 144 347 160 381
rect 194 347 210 381
rect 144 331 210 347
rect 262 381 328 397
rect 262 347 278 381
rect 312 347 328 381
rect 262 331 328 347
rect 380 381 446 397
rect 380 347 396 381
rect 430 347 446 381
rect 380 331 446 347
rect 498 381 564 397
rect 498 347 514 381
rect 548 347 564 381
rect 498 331 564 347
rect -561 300 -501 331
rect -443 300 -383 331
rect -325 300 -265 331
rect -207 300 -147 331
rect -89 300 -29 331
rect 29 300 89 331
rect 147 300 207 331
rect 265 300 325 331
rect 383 300 443 331
rect 501 300 561 331
rect -561 -331 -501 -300
rect -443 -331 -383 -300
rect -325 -331 -265 -300
rect -207 -331 -147 -300
rect -89 -331 -29 -300
rect 29 -331 89 -300
rect 147 -331 207 -300
rect 265 -331 325 -300
rect 383 -331 443 -300
rect 501 -331 561 -300
rect -564 -347 -498 -331
rect -564 -381 -548 -347
rect -514 -381 -498 -347
rect -564 -397 -498 -381
rect -446 -347 -380 -331
rect -446 -381 -430 -347
rect -396 -381 -380 -347
rect -446 -397 -380 -381
rect -328 -347 -262 -331
rect -328 -381 -312 -347
rect -278 -381 -262 -347
rect -328 -397 -262 -381
rect -210 -347 -144 -331
rect -210 -381 -194 -347
rect -160 -381 -144 -347
rect -210 -397 -144 -381
rect -92 -347 -26 -331
rect -92 -381 -76 -347
rect -42 -381 -26 -347
rect -92 -397 -26 -381
rect 26 -347 92 -331
rect 26 -381 42 -347
rect 76 -381 92 -347
rect 26 -397 92 -381
rect 144 -347 210 -331
rect 144 -381 160 -347
rect 194 -381 210 -347
rect 144 -397 210 -381
rect 262 -347 328 -331
rect 262 -381 278 -347
rect 312 -381 328 -347
rect 262 -397 328 -381
rect 380 -347 446 -331
rect 380 -381 396 -347
rect 430 -381 446 -347
rect 380 -397 446 -381
rect 498 -347 564 -331
rect 498 -381 514 -347
rect 548 -381 564 -347
rect 498 -397 564 -381
rect -564 -455 -498 -439
rect -564 -489 -548 -455
rect -514 -489 -498 -455
rect -564 -505 -498 -489
rect -446 -455 -380 -439
rect -446 -489 -430 -455
rect -396 -489 -380 -455
rect -446 -505 -380 -489
rect -328 -455 -262 -439
rect -328 -489 -312 -455
rect -278 -489 -262 -455
rect -328 -505 -262 -489
rect -210 -455 -144 -439
rect -210 -489 -194 -455
rect -160 -489 -144 -455
rect -210 -505 -144 -489
rect -92 -455 -26 -439
rect -92 -489 -76 -455
rect -42 -489 -26 -455
rect -92 -505 -26 -489
rect 26 -455 92 -439
rect 26 -489 42 -455
rect 76 -489 92 -455
rect 26 -505 92 -489
rect 144 -455 210 -439
rect 144 -489 160 -455
rect 194 -489 210 -455
rect 144 -505 210 -489
rect 262 -455 328 -439
rect 262 -489 278 -455
rect 312 -489 328 -455
rect 262 -505 328 -489
rect 380 -455 446 -439
rect 380 -489 396 -455
rect 430 -489 446 -455
rect 380 -505 446 -489
rect 498 -455 564 -439
rect 498 -489 514 -455
rect 548 -489 564 -455
rect 498 -505 564 -489
rect -561 -536 -501 -505
rect -443 -536 -383 -505
rect -325 -536 -265 -505
rect -207 -536 -147 -505
rect -89 -536 -29 -505
rect 29 -536 89 -505
rect 147 -536 207 -505
rect 265 -536 325 -505
rect 383 -536 443 -505
rect 501 -536 561 -505
rect -561 -1167 -501 -1136
rect -443 -1167 -383 -1136
rect -325 -1167 -265 -1136
rect -207 -1167 -147 -1136
rect -89 -1167 -29 -1136
rect 29 -1167 89 -1136
rect 147 -1167 207 -1136
rect 265 -1167 325 -1136
rect 383 -1167 443 -1136
rect 501 -1167 561 -1136
rect -564 -1183 -498 -1167
rect -564 -1217 -548 -1183
rect -514 -1217 -498 -1183
rect -564 -1233 -498 -1217
rect -446 -1183 -380 -1167
rect -446 -1217 -430 -1183
rect -396 -1217 -380 -1183
rect -446 -1233 -380 -1217
rect -328 -1183 -262 -1167
rect -328 -1217 -312 -1183
rect -278 -1217 -262 -1183
rect -328 -1233 -262 -1217
rect -210 -1183 -144 -1167
rect -210 -1217 -194 -1183
rect -160 -1217 -144 -1183
rect -210 -1233 -144 -1217
rect -92 -1183 -26 -1167
rect -92 -1217 -76 -1183
rect -42 -1217 -26 -1183
rect -92 -1233 -26 -1217
rect 26 -1183 92 -1167
rect 26 -1217 42 -1183
rect 76 -1217 92 -1183
rect 26 -1233 92 -1217
rect 144 -1183 210 -1167
rect 144 -1217 160 -1183
rect 194 -1217 210 -1183
rect 144 -1233 210 -1217
rect 262 -1183 328 -1167
rect 262 -1217 278 -1183
rect 312 -1217 328 -1183
rect 262 -1233 328 -1217
rect 380 -1183 446 -1167
rect 380 -1217 396 -1183
rect 430 -1217 446 -1183
rect 380 -1233 446 -1217
rect 498 -1183 564 -1167
rect 498 -1217 514 -1183
rect 548 -1217 564 -1183
rect 498 -1233 564 -1217
<< polycont >>
rect -548 1183 -514 1217
rect -430 1183 -396 1217
rect -312 1183 -278 1217
rect -194 1183 -160 1217
rect -76 1183 -42 1217
rect 42 1183 76 1217
rect 160 1183 194 1217
rect 278 1183 312 1217
rect 396 1183 430 1217
rect 514 1183 548 1217
rect -548 455 -514 489
rect -430 455 -396 489
rect -312 455 -278 489
rect -194 455 -160 489
rect -76 455 -42 489
rect 42 455 76 489
rect 160 455 194 489
rect 278 455 312 489
rect 396 455 430 489
rect 514 455 548 489
rect -548 347 -514 381
rect -430 347 -396 381
rect -312 347 -278 381
rect -194 347 -160 381
rect -76 347 -42 381
rect 42 347 76 381
rect 160 347 194 381
rect 278 347 312 381
rect 396 347 430 381
rect 514 347 548 381
rect -548 -381 -514 -347
rect -430 -381 -396 -347
rect -312 -381 -278 -347
rect -194 -381 -160 -347
rect -76 -381 -42 -347
rect 42 -381 76 -347
rect 160 -381 194 -347
rect 278 -381 312 -347
rect 396 -381 430 -347
rect 514 -381 548 -347
rect -548 -489 -514 -455
rect -430 -489 -396 -455
rect -312 -489 -278 -455
rect -194 -489 -160 -455
rect -76 -489 -42 -455
rect 42 -489 76 -455
rect 160 -489 194 -455
rect 278 -489 312 -455
rect 396 -489 430 -455
rect 514 -489 548 -455
rect -548 -1217 -514 -1183
rect -430 -1217 -396 -1183
rect -312 -1217 -278 -1183
rect -194 -1217 -160 -1183
rect -76 -1217 -42 -1183
rect 42 -1217 76 -1183
rect 160 -1217 194 -1183
rect 278 -1217 312 -1183
rect 396 -1217 430 -1183
rect 514 -1217 548 -1183
<< locali >>
rect -721 1285 -625 1319
rect 625 1285 721 1319
rect -721 1223 -687 1285
rect 687 1223 721 1285
rect -564 1183 -548 1217
rect -514 1183 -498 1217
rect -446 1183 -430 1217
rect -396 1183 -380 1217
rect -328 1183 -312 1217
rect -278 1183 -262 1217
rect -210 1183 -194 1217
rect -160 1183 -144 1217
rect -92 1183 -76 1217
rect -42 1183 -26 1217
rect 26 1183 42 1217
rect 76 1183 92 1217
rect 144 1183 160 1217
rect 194 1183 210 1217
rect 262 1183 278 1217
rect 312 1183 328 1217
rect 380 1183 396 1217
rect 430 1183 446 1217
rect 498 1183 514 1217
rect 548 1183 564 1217
rect -607 1124 -573 1140
rect -607 532 -573 548
rect -489 1124 -455 1140
rect -489 532 -455 548
rect -371 1124 -337 1140
rect -371 532 -337 548
rect -253 1124 -219 1140
rect -253 532 -219 548
rect -135 1124 -101 1140
rect -135 532 -101 548
rect -17 1124 17 1140
rect -17 532 17 548
rect 101 1124 135 1140
rect 101 532 135 548
rect 219 1124 253 1140
rect 219 532 253 548
rect 337 1124 371 1140
rect 337 532 371 548
rect 455 1124 489 1140
rect 455 532 489 548
rect 573 1124 607 1140
rect 573 532 607 548
rect -564 455 -548 489
rect -514 455 -498 489
rect -446 455 -430 489
rect -396 455 -380 489
rect -328 455 -312 489
rect -278 455 -262 489
rect -210 455 -194 489
rect -160 455 -144 489
rect -92 455 -76 489
rect -42 455 -26 489
rect 26 455 42 489
rect 76 455 92 489
rect 144 455 160 489
rect 194 455 210 489
rect 262 455 278 489
rect 312 455 328 489
rect 380 455 396 489
rect 430 455 446 489
rect 498 455 514 489
rect 548 455 564 489
rect -564 347 -548 381
rect -514 347 -498 381
rect -446 347 -430 381
rect -396 347 -380 381
rect -328 347 -312 381
rect -278 347 -262 381
rect -210 347 -194 381
rect -160 347 -144 381
rect -92 347 -76 381
rect -42 347 -26 381
rect 26 347 42 381
rect 76 347 92 381
rect 144 347 160 381
rect 194 347 210 381
rect 262 347 278 381
rect 312 347 328 381
rect 380 347 396 381
rect 430 347 446 381
rect 498 347 514 381
rect 548 347 564 381
rect -607 288 -573 304
rect -607 -304 -573 -288
rect -489 288 -455 304
rect -489 -304 -455 -288
rect -371 288 -337 304
rect -371 -304 -337 -288
rect -253 288 -219 304
rect -253 -304 -219 -288
rect -135 288 -101 304
rect -135 -304 -101 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 101 288 135 304
rect 101 -304 135 -288
rect 219 288 253 304
rect 219 -304 253 -288
rect 337 288 371 304
rect 337 -304 371 -288
rect 455 288 489 304
rect 455 -304 489 -288
rect 573 288 607 304
rect 573 -304 607 -288
rect -564 -381 -548 -347
rect -514 -381 -498 -347
rect -446 -381 -430 -347
rect -396 -381 -380 -347
rect -328 -381 -312 -347
rect -278 -381 -262 -347
rect -210 -381 -194 -347
rect -160 -381 -144 -347
rect -92 -381 -76 -347
rect -42 -381 -26 -347
rect 26 -381 42 -347
rect 76 -381 92 -347
rect 144 -381 160 -347
rect 194 -381 210 -347
rect 262 -381 278 -347
rect 312 -381 328 -347
rect 380 -381 396 -347
rect 430 -381 446 -347
rect 498 -381 514 -347
rect 548 -381 564 -347
rect -564 -489 -548 -455
rect -514 -489 -498 -455
rect -446 -489 -430 -455
rect -396 -489 -380 -455
rect -328 -489 -312 -455
rect -278 -489 -262 -455
rect -210 -489 -194 -455
rect -160 -489 -144 -455
rect -92 -489 -76 -455
rect -42 -489 -26 -455
rect 26 -489 42 -455
rect 76 -489 92 -455
rect 144 -489 160 -455
rect 194 -489 210 -455
rect 262 -489 278 -455
rect 312 -489 328 -455
rect 380 -489 396 -455
rect 430 -489 446 -455
rect 498 -489 514 -455
rect 548 -489 564 -455
rect -607 -548 -573 -532
rect -607 -1140 -573 -1124
rect -489 -548 -455 -532
rect -489 -1140 -455 -1124
rect -371 -548 -337 -532
rect -371 -1140 -337 -1124
rect -253 -548 -219 -532
rect -253 -1140 -219 -1124
rect -135 -548 -101 -532
rect -135 -1140 -101 -1124
rect -17 -548 17 -532
rect -17 -1140 17 -1124
rect 101 -548 135 -532
rect 101 -1140 135 -1124
rect 219 -548 253 -532
rect 219 -1140 253 -1124
rect 337 -548 371 -532
rect 337 -1140 371 -1124
rect 455 -548 489 -532
rect 455 -1140 489 -1124
rect 573 -548 607 -532
rect 573 -1140 607 -1124
rect -564 -1217 -548 -1183
rect -514 -1217 -498 -1183
rect -446 -1217 -430 -1183
rect -396 -1217 -380 -1183
rect -328 -1217 -312 -1183
rect -278 -1217 -262 -1183
rect -210 -1217 -194 -1183
rect -160 -1217 -144 -1183
rect -92 -1217 -76 -1183
rect -42 -1217 -26 -1183
rect 26 -1217 42 -1183
rect 76 -1217 92 -1183
rect 144 -1217 160 -1183
rect 194 -1217 210 -1183
rect 262 -1217 278 -1183
rect 312 -1217 328 -1183
rect 380 -1217 396 -1183
rect 430 -1217 446 -1183
rect 498 -1217 514 -1183
rect 548 -1217 564 -1183
rect -721 -1285 -687 -1223
rect 687 -1285 721 -1223
rect -721 -1319 -625 -1285
rect 625 -1319 721 -1285
<< viali >>
rect -548 1183 -514 1217
rect -430 1183 -396 1217
rect -312 1183 -278 1217
rect -194 1183 -160 1217
rect -76 1183 -42 1217
rect 42 1183 76 1217
rect 160 1183 194 1217
rect 278 1183 312 1217
rect 396 1183 430 1217
rect 514 1183 548 1217
rect -607 548 -573 1124
rect -489 548 -455 1124
rect -371 548 -337 1124
rect -253 548 -219 1124
rect -135 548 -101 1124
rect -17 548 17 1124
rect 101 548 135 1124
rect 219 548 253 1124
rect 337 548 371 1124
rect 455 548 489 1124
rect 573 548 607 1124
rect -548 455 -514 489
rect -430 455 -396 489
rect -312 455 -278 489
rect -194 455 -160 489
rect -76 455 -42 489
rect 42 455 76 489
rect 160 455 194 489
rect 278 455 312 489
rect 396 455 430 489
rect 514 455 548 489
rect -548 347 -514 381
rect -430 347 -396 381
rect -312 347 -278 381
rect -194 347 -160 381
rect -76 347 -42 381
rect 42 347 76 381
rect 160 347 194 381
rect 278 347 312 381
rect 396 347 430 381
rect 514 347 548 381
rect -607 -288 -573 288
rect -489 -288 -455 288
rect -371 -288 -337 288
rect -253 -288 -219 288
rect -135 -288 -101 288
rect -17 -288 17 288
rect 101 -288 135 288
rect 219 -288 253 288
rect 337 -288 371 288
rect 455 -288 489 288
rect 573 -288 607 288
rect -548 -381 -514 -347
rect -430 -381 -396 -347
rect -312 -381 -278 -347
rect -194 -381 -160 -347
rect -76 -381 -42 -347
rect 42 -381 76 -347
rect 160 -381 194 -347
rect 278 -381 312 -347
rect 396 -381 430 -347
rect 514 -381 548 -347
rect -548 -489 -514 -455
rect -430 -489 -396 -455
rect -312 -489 -278 -455
rect -194 -489 -160 -455
rect -76 -489 -42 -455
rect 42 -489 76 -455
rect 160 -489 194 -455
rect 278 -489 312 -455
rect 396 -489 430 -455
rect 514 -489 548 -455
rect -607 -1124 -573 -548
rect -489 -1124 -455 -548
rect -371 -1124 -337 -548
rect -253 -1124 -219 -548
rect -135 -1124 -101 -548
rect -17 -1124 17 -548
rect 101 -1124 135 -548
rect 219 -1124 253 -548
rect 337 -1124 371 -548
rect 455 -1124 489 -548
rect 573 -1124 607 -548
rect -548 -1217 -514 -1183
rect -430 -1217 -396 -1183
rect -312 -1217 -278 -1183
rect -194 -1217 -160 -1183
rect -76 -1217 -42 -1183
rect 42 -1217 76 -1183
rect 160 -1217 194 -1183
rect 278 -1217 312 -1183
rect 396 -1217 430 -1183
rect 514 -1217 548 -1183
<< metal1 >>
rect -560 1217 -502 1223
rect -560 1183 -548 1217
rect -514 1183 -502 1217
rect -560 1177 -502 1183
rect -442 1217 -384 1223
rect -442 1183 -430 1217
rect -396 1183 -384 1217
rect -442 1177 -384 1183
rect -324 1217 -266 1223
rect -324 1183 -312 1217
rect -278 1183 -266 1217
rect -324 1177 -266 1183
rect -206 1217 -148 1223
rect -206 1183 -194 1217
rect -160 1183 -148 1217
rect -206 1177 -148 1183
rect -88 1217 -30 1223
rect -88 1183 -76 1217
rect -42 1183 -30 1217
rect -88 1177 -30 1183
rect 30 1217 88 1223
rect 30 1183 42 1217
rect 76 1183 88 1217
rect 30 1177 88 1183
rect 148 1217 206 1223
rect 148 1183 160 1217
rect 194 1183 206 1217
rect 148 1177 206 1183
rect 266 1217 324 1223
rect 266 1183 278 1217
rect 312 1183 324 1217
rect 266 1177 324 1183
rect 384 1217 442 1223
rect 384 1183 396 1217
rect 430 1183 442 1217
rect 384 1177 442 1183
rect 502 1217 560 1223
rect 502 1183 514 1217
rect 548 1183 560 1217
rect 502 1177 560 1183
rect -613 1124 -567 1136
rect -613 548 -607 1124
rect -573 548 -567 1124
rect -613 536 -567 548
rect -495 1124 -449 1136
rect -495 548 -489 1124
rect -455 548 -449 1124
rect -495 536 -449 548
rect -377 1124 -331 1136
rect -377 548 -371 1124
rect -337 548 -331 1124
rect -377 536 -331 548
rect -259 1124 -213 1136
rect -259 548 -253 1124
rect -219 548 -213 1124
rect -259 536 -213 548
rect -141 1124 -95 1136
rect -141 548 -135 1124
rect -101 548 -95 1124
rect -141 536 -95 548
rect -23 1124 23 1136
rect -23 548 -17 1124
rect 17 548 23 1124
rect -23 536 23 548
rect 95 1124 141 1136
rect 95 548 101 1124
rect 135 548 141 1124
rect 95 536 141 548
rect 213 1124 259 1136
rect 213 548 219 1124
rect 253 548 259 1124
rect 213 536 259 548
rect 331 1124 377 1136
rect 331 548 337 1124
rect 371 548 377 1124
rect 331 536 377 548
rect 449 1124 495 1136
rect 449 548 455 1124
rect 489 548 495 1124
rect 449 536 495 548
rect 567 1124 613 1136
rect 567 548 573 1124
rect 607 548 613 1124
rect 567 536 613 548
rect -560 489 -502 495
rect -560 455 -548 489
rect -514 455 -502 489
rect -560 449 -502 455
rect -442 489 -384 495
rect -442 455 -430 489
rect -396 455 -384 489
rect -442 449 -384 455
rect -324 489 -266 495
rect -324 455 -312 489
rect -278 455 -266 489
rect -324 449 -266 455
rect -206 489 -148 495
rect -206 455 -194 489
rect -160 455 -148 489
rect -206 449 -148 455
rect -88 489 -30 495
rect -88 455 -76 489
rect -42 455 -30 489
rect -88 449 -30 455
rect 30 489 88 495
rect 30 455 42 489
rect 76 455 88 489
rect 30 449 88 455
rect 148 489 206 495
rect 148 455 160 489
rect 194 455 206 489
rect 148 449 206 455
rect 266 489 324 495
rect 266 455 278 489
rect 312 455 324 489
rect 266 449 324 455
rect 384 489 442 495
rect 384 455 396 489
rect 430 455 442 489
rect 384 449 442 455
rect 502 489 560 495
rect 502 455 514 489
rect 548 455 560 489
rect 502 449 560 455
rect -560 381 -502 387
rect -560 347 -548 381
rect -514 347 -502 381
rect -560 341 -502 347
rect -442 381 -384 387
rect -442 347 -430 381
rect -396 347 -384 381
rect -442 341 -384 347
rect -324 381 -266 387
rect -324 347 -312 381
rect -278 347 -266 381
rect -324 341 -266 347
rect -206 381 -148 387
rect -206 347 -194 381
rect -160 347 -148 381
rect -206 341 -148 347
rect -88 381 -30 387
rect -88 347 -76 381
rect -42 347 -30 381
rect -88 341 -30 347
rect 30 381 88 387
rect 30 347 42 381
rect 76 347 88 381
rect 30 341 88 347
rect 148 381 206 387
rect 148 347 160 381
rect 194 347 206 381
rect 148 341 206 347
rect 266 381 324 387
rect 266 347 278 381
rect 312 347 324 381
rect 266 341 324 347
rect 384 381 442 387
rect 384 347 396 381
rect 430 347 442 381
rect 384 341 442 347
rect 502 381 560 387
rect 502 347 514 381
rect 548 347 560 381
rect 502 341 560 347
rect -613 288 -567 300
rect -613 -288 -607 288
rect -573 -288 -567 288
rect -613 -300 -567 -288
rect -495 288 -449 300
rect -495 -288 -489 288
rect -455 -288 -449 288
rect -495 -300 -449 -288
rect -377 288 -331 300
rect -377 -288 -371 288
rect -337 -288 -331 288
rect -377 -300 -331 -288
rect -259 288 -213 300
rect -259 -288 -253 288
rect -219 -288 -213 288
rect -259 -300 -213 -288
rect -141 288 -95 300
rect -141 -288 -135 288
rect -101 -288 -95 288
rect -141 -300 -95 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 95 288 141 300
rect 95 -288 101 288
rect 135 -288 141 288
rect 95 -300 141 -288
rect 213 288 259 300
rect 213 -288 219 288
rect 253 -288 259 288
rect 213 -300 259 -288
rect 331 288 377 300
rect 331 -288 337 288
rect 371 -288 377 288
rect 331 -300 377 -288
rect 449 288 495 300
rect 449 -288 455 288
rect 489 -288 495 288
rect 449 -300 495 -288
rect 567 288 613 300
rect 567 -288 573 288
rect 607 -288 613 288
rect 567 -300 613 -288
rect -560 -347 -502 -341
rect -560 -381 -548 -347
rect -514 -381 -502 -347
rect -560 -387 -502 -381
rect -442 -347 -384 -341
rect -442 -381 -430 -347
rect -396 -381 -384 -347
rect -442 -387 -384 -381
rect -324 -347 -266 -341
rect -324 -381 -312 -347
rect -278 -381 -266 -347
rect -324 -387 -266 -381
rect -206 -347 -148 -341
rect -206 -381 -194 -347
rect -160 -381 -148 -347
rect -206 -387 -148 -381
rect -88 -347 -30 -341
rect -88 -381 -76 -347
rect -42 -381 -30 -347
rect -88 -387 -30 -381
rect 30 -347 88 -341
rect 30 -381 42 -347
rect 76 -381 88 -347
rect 30 -387 88 -381
rect 148 -347 206 -341
rect 148 -381 160 -347
rect 194 -381 206 -347
rect 148 -387 206 -381
rect 266 -347 324 -341
rect 266 -381 278 -347
rect 312 -381 324 -347
rect 266 -387 324 -381
rect 384 -347 442 -341
rect 384 -381 396 -347
rect 430 -381 442 -347
rect 384 -387 442 -381
rect 502 -347 560 -341
rect 502 -381 514 -347
rect 548 -381 560 -347
rect 502 -387 560 -381
rect -560 -455 -502 -449
rect -560 -489 -548 -455
rect -514 -489 -502 -455
rect -560 -495 -502 -489
rect -442 -455 -384 -449
rect -442 -489 -430 -455
rect -396 -489 -384 -455
rect -442 -495 -384 -489
rect -324 -455 -266 -449
rect -324 -489 -312 -455
rect -278 -489 -266 -455
rect -324 -495 -266 -489
rect -206 -455 -148 -449
rect -206 -489 -194 -455
rect -160 -489 -148 -455
rect -206 -495 -148 -489
rect -88 -455 -30 -449
rect -88 -489 -76 -455
rect -42 -489 -30 -455
rect -88 -495 -30 -489
rect 30 -455 88 -449
rect 30 -489 42 -455
rect 76 -489 88 -455
rect 30 -495 88 -489
rect 148 -455 206 -449
rect 148 -489 160 -455
rect 194 -489 206 -455
rect 148 -495 206 -489
rect 266 -455 324 -449
rect 266 -489 278 -455
rect 312 -489 324 -455
rect 266 -495 324 -489
rect 384 -455 442 -449
rect 384 -489 396 -455
rect 430 -489 442 -455
rect 384 -495 442 -489
rect 502 -455 560 -449
rect 502 -489 514 -455
rect 548 -489 560 -455
rect 502 -495 560 -489
rect -613 -548 -567 -536
rect -613 -1124 -607 -548
rect -573 -1124 -567 -548
rect -613 -1136 -567 -1124
rect -495 -548 -449 -536
rect -495 -1124 -489 -548
rect -455 -1124 -449 -548
rect -495 -1136 -449 -1124
rect -377 -548 -331 -536
rect -377 -1124 -371 -548
rect -337 -1124 -331 -548
rect -377 -1136 -331 -1124
rect -259 -548 -213 -536
rect -259 -1124 -253 -548
rect -219 -1124 -213 -548
rect -259 -1136 -213 -1124
rect -141 -548 -95 -536
rect -141 -1124 -135 -548
rect -101 -1124 -95 -548
rect -141 -1136 -95 -1124
rect -23 -548 23 -536
rect -23 -1124 -17 -548
rect 17 -1124 23 -548
rect -23 -1136 23 -1124
rect 95 -548 141 -536
rect 95 -1124 101 -548
rect 135 -1124 141 -548
rect 95 -1136 141 -1124
rect 213 -548 259 -536
rect 213 -1124 219 -548
rect 253 -1124 259 -548
rect 213 -1136 259 -1124
rect 331 -548 377 -536
rect 331 -1124 337 -548
rect 371 -1124 377 -548
rect 331 -1136 377 -1124
rect 449 -548 495 -536
rect 449 -1124 455 -548
rect 489 -1124 495 -548
rect 449 -1136 495 -1124
rect 567 -548 613 -536
rect 567 -1124 573 -548
rect 607 -1124 613 -548
rect 567 -1136 613 -1124
rect -560 -1183 -502 -1177
rect -560 -1217 -548 -1183
rect -514 -1217 -502 -1183
rect -560 -1223 -502 -1217
rect -442 -1183 -384 -1177
rect -442 -1217 -430 -1183
rect -396 -1217 -384 -1183
rect -442 -1223 -384 -1217
rect -324 -1183 -266 -1177
rect -324 -1217 -312 -1183
rect -278 -1217 -266 -1183
rect -324 -1223 -266 -1217
rect -206 -1183 -148 -1177
rect -206 -1217 -194 -1183
rect -160 -1217 -148 -1183
rect -206 -1223 -148 -1217
rect -88 -1183 -30 -1177
rect -88 -1217 -76 -1183
rect -42 -1217 -30 -1183
rect -88 -1223 -30 -1217
rect 30 -1183 88 -1177
rect 30 -1217 42 -1183
rect 76 -1217 88 -1183
rect 30 -1223 88 -1217
rect 148 -1183 206 -1177
rect 148 -1217 160 -1183
rect 194 -1217 206 -1183
rect 148 -1223 206 -1217
rect 266 -1183 324 -1177
rect 266 -1217 278 -1183
rect 312 -1217 324 -1183
rect 266 -1223 324 -1217
rect 384 -1183 442 -1177
rect 384 -1217 396 -1183
rect 430 -1217 442 -1183
rect 384 -1223 442 -1217
rect 502 -1183 560 -1177
rect 502 -1217 514 -1183
rect 548 -1217 560 -1183
rect 502 -1223 560 -1217
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -704 -1302 704 1302
string parameters w 3 l 0.3 m 3 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
