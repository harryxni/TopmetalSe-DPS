magic
tech sky130B
magscale 1 2
timestamp 1606424956
<< metal3 >>
rect -1686 1572 1686 1600
rect -1686 -1572 1602 1572
rect 1666 -1572 1686 1572
rect -1686 -1600 1686 -1572
<< via3 >>
rect 1602 -1572 1666 1572
<< mimcap >>
rect -1586 1460 1414 1500
rect -1586 -1460 -1546 1460
rect 1374 -1460 1414 1460
rect -1586 -1500 1414 -1460
<< mimcapcontact >>
rect -1546 -1460 1374 1460
<< metal4 >>
rect 1586 1572 1682 1588
rect -1547 1460 1375 1461
rect -1547 -1460 -1546 1460
rect 1374 -1460 1375 1460
rect -1547 -1461 1375 -1460
rect 1586 -1572 1602 1572
rect 1666 -1572 1682 1572
rect 1586 -1588 1682 -1572
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -1686 -1600 1514 1600
string parameters w 15 l 15 val 235.2 carea 1.00 cperi 0.17 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1
string library sky130
<< end >>
