magic
tech sky130B
magscale 1 2
timestamp 1607649912
<< nwell >>
rect -8177 -1537 8177 1537
<< pmos >>
rect -7981 118 -7861 1318
rect -7803 118 -7683 1318
rect -7625 118 -7505 1318
rect -7447 118 -7327 1318
rect -7269 118 -7149 1318
rect -7091 118 -6971 1318
rect -6913 118 -6793 1318
rect -6735 118 -6615 1318
rect -6557 118 -6437 1318
rect -6379 118 -6259 1318
rect -6201 118 -6081 1318
rect -6023 118 -5903 1318
rect -5845 118 -5725 1318
rect -5667 118 -5547 1318
rect -5489 118 -5369 1318
rect -5311 118 -5191 1318
rect -5133 118 -5013 1318
rect -4955 118 -4835 1318
rect -4777 118 -4657 1318
rect -4599 118 -4479 1318
rect -4421 118 -4301 1318
rect -4243 118 -4123 1318
rect -4065 118 -3945 1318
rect -3887 118 -3767 1318
rect -3709 118 -3589 1318
rect -3531 118 -3411 1318
rect -3353 118 -3233 1318
rect -3175 118 -3055 1318
rect -2997 118 -2877 1318
rect -2819 118 -2699 1318
rect -2641 118 -2521 1318
rect -2463 118 -2343 1318
rect -2285 118 -2165 1318
rect -2107 118 -1987 1318
rect -1929 118 -1809 1318
rect -1751 118 -1631 1318
rect -1573 118 -1453 1318
rect -1395 118 -1275 1318
rect -1217 118 -1097 1318
rect -1039 118 -919 1318
rect -861 118 -741 1318
rect -683 118 -563 1318
rect -505 118 -385 1318
rect -327 118 -207 1318
rect -149 118 -29 1318
rect 29 118 149 1318
rect 207 118 327 1318
rect 385 118 505 1318
rect 563 118 683 1318
rect 741 118 861 1318
rect 919 118 1039 1318
rect 1097 118 1217 1318
rect 1275 118 1395 1318
rect 1453 118 1573 1318
rect 1631 118 1751 1318
rect 1809 118 1929 1318
rect 1987 118 2107 1318
rect 2165 118 2285 1318
rect 2343 118 2463 1318
rect 2521 118 2641 1318
rect 2699 118 2819 1318
rect 2877 118 2997 1318
rect 3055 118 3175 1318
rect 3233 118 3353 1318
rect 3411 118 3531 1318
rect 3589 118 3709 1318
rect 3767 118 3887 1318
rect 3945 118 4065 1318
rect 4123 118 4243 1318
rect 4301 118 4421 1318
rect 4479 118 4599 1318
rect 4657 118 4777 1318
rect 4835 118 4955 1318
rect 5013 118 5133 1318
rect 5191 118 5311 1318
rect 5369 118 5489 1318
rect 5547 118 5667 1318
rect 5725 118 5845 1318
rect 5903 118 6023 1318
rect 6081 118 6201 1318
rect 6259 118 6379 1318
rect 6437 118 6557 1318
rect 6615 118 6735 1318
rect 6793 118 6913 1318
rect 6971 118 7091 1318
rect 7149 118 7269 1318
rect 7327 118 7447 1318
rect 7505 118 7625 1318
rect 7683 118 7803 1318
rect 7861 118 7981 1318
rect -7981 -1318 -7861 -118
rect -7803 -1318 -7683 -118
rect -7625 -1318 -7505 -118
rect -7447 -1318 -7327 -118
rect -7269 -1318 -7149 -118
rect -7091 -1318 -6971 -118
rect -6913 -1318 -6793 -118
rect -6735 -1318 -6615 -118
rect -6557 -1318 -6437 -118
rect -6379 -1318 -6259 -118
rect -6201 -1318 -6081 -118
rect -6023 -1318 -5903 -118
rect -5845 -1318 -5725 -118
rect -5667 -1318 -5547 -118
rect -5489 -1318 -5369 -118
rect -5311 -1318 -5191 -118
rect -5133 -1318 -5013 -118
rect -4955 -1318 -4835 -118
rect -4777 -1318 -4657 -118
rect -4599 -1318 -4479 -118
rect -4421 -1318 -4301 -118
rect -4243 -1318 -4123 -118
rect -4065 -1318 -3945 -118
rect -3887 -1318 -3767 -118
rect -3709 -1318 -3589 -118
rect -3531 -1318 -3411 -118
rect -3353 -1318 -3233 -118
rect -3175 -1318 -3055 -118
rect -2997 -1318 -2877 -118
rect -2819 -1318 -2699 -118
rect -2641 -1318 -2521 -118
rect -2463 -1318 -2343 -118
rect -2285 -1318 -2165 -118
rect -2107 -1318 -1987 -118
rect -1929 -1318 -1809 -118
rect -1751 -1318 -1631 -118
rect -1573 -1318 -1453 -118
rect -1395 -1318 -1275 -118
rect -1217 -1318 -1097 -118
rect -1039 -1318 -919 -118
rect -861 -1318 -741 -118
rect -683 -1318 -563 -118
rect -505 -1318 -385 -118
rect -327 -1318 -207 -118
rect -149 -1318 -29 -118
rect 29 -1318 149 -118
rect 207 -1318 327 -118
rect 385 -1318 505 -118
rect 563 -1318 683 -118
rect 741 -1318 861 -118
rect 919 -1318 1039 -118
rect 1097 -1318 1217 -118
rect 1275 -1318 1395 -118
rect 1453 -1318 1573 -118
rect 1631 -1318 1751 -118
rect 1809 -1318 1929 -118
rect 1987 -1318 2107 -118
rect 2165 -1318 2285 -118
rect 2343 -1318 2463 -118
rect 2521 -1318 2641 -118
rect 2699 -1318 2819 -118
rect 2877 -1318 2997 -118
rect 3055 -1318 3175 -118
rect 3233 -1318 3353 -118
rect 3411 -1318 3531 -118
rect 3589 -1318 3709 -118
rect 3767 -1318 3887 -118
rect 3945 -1318 4065 -118
rect 4123 -1318 4243 -118
rect 4301 -1318 4421 -118
rect 4479 -1318 4599 -118
rect 4657 -1318 4777 -118
rect 4835 -1318 4955 -118
rect 5013 -1318 5133 -118
rect 5191 -1318 5311 -118
rect 5369 -1318 5489 -118
rect 5547 -1318 5667 -118
rect 5725 -1318 5845 -118
rect 5903 -1318 6023 -118
rect 6081 -1318 6201 -118
rect 6259 -1318 6379 -118
rect 6437 -1318 6557 -118
rect 6615 -1318 6735 -118
rect 6793 -1318 6913 -118
rect 6971 -1318 7091 -118
rect 7149 -1318 7269 -118
rect 7327 -1318 7447 -118
rect 7505 -1318 7625 -118
rect 7683 -1318 7803 -118
rect 7861 -1318 7981 -118
<< pdiff >>
rect -8039 1306 -7981 1318
rect -8039 130 -8027 1306
rect -7993 130 -7981 1306
rect -8039 118 -7981 130
rect -7861 1306 -7803 1318
rect -7861 130 -7849 1306
rect -7815 130 -7803 1306
rect -7861 118 -7803 130
rect -7683 1306 -7625 1318
rect -7683 130 -7671 1306
rect -7637 130 -7625 1306
rect -7683 118 -7625 130
rect -7505 1306 -7447 1318
rect -7505 130 -7493 1306
rect -7459 130 -7447 1306
rect -7505 118 -7447 130
rect -7327 1306 -7269 1318
rect -7327 130 -7315 1306
rect -7281 130 -7269 1306
rect -7327 118 -7269 130
rect -7149 1306 -7091 1318
rect -7149 130 -7137 1306
rect -7103 130 -7091 1306
rect -7149 118 -7091 130
rect -6971 1306 -6913 1318
rect -6971 130 -6959 1306
rect -6925 130 -6913 1306
rect -6971 118 -6913 130
rect -6793 1306 -6735 1318
rect -6793 130 -6781 1306
rect -6747 130 -6735 1306
rect -6793 118 -6735 130
rect -6615 1306 -6557 1318
rect -6615 130 -6603 1306
rect -6569 130 -6557 1306
rect -6615 118 -6557 130
rect -6437 1306 -6379 1318
rect -6437 130 -6425 1306
rect -6391 130 -6379 1306
rect -6437 118 -6379 130
rect -6259 1306 -6201 1318
rect -6259 130 -6247 1306
rect -6213 130 -6201 1306
rect -6259 118 -6201 130
rect -6081 1306 -6023 1318
rect -6081 130 -6069 1306
rect -6035 130 -6023 1306
rect -6081 118 -6023 130
rect -5903 1306 -5845 1318
rect -5903 130 -5891 1306
rect -5857 130 -5845 1306
rect -5903 118 -5845 130
rect -5725 1306 -5667 1318
rect -5725 130 -5713 1306
rect -5679 130 -5667 1306
rect -5725 118 -5667 130
rect -5547 1306 -5489 1318
rect -5547 130 -5535 1306
rect -5501 130 -5489 1306
rect -5547 118 -5489 130
rect -5369 1306 -5311 1318
rect -5369 130 -5357 1306
rect -5323 130 -5311 1306
rect -5369 118 -5311 130
rect -5191 1306 -5133 1318
rect -5191 130 -5179 1306
rect -5145 130 -5133 1306
rect -5191 118 -5133 130
rect -5013 1306 -4955 1318
rect -5013 130 -5001 1306
rect -4967 130 -4955 1306
rect -5013 118 -4955 130
rect -4835 1306 -4777 1318
rect -4835 130 -4823 1306
rect -4789 130 -4777 1306
rect -4835 118 -4777 130
rect -4657 1306 -4599 1318
rect -4657 130 -4645 1306
rect -4611 130 -4599 1306
rect -4657 118 -4599 130
rect -4479 1306 -4421 1318
rect -4479 130 -4467 1306
rect -4433 130 -4421 1306
rect -4479 118 -4421 130
rect -4301 1306 -4243 1318
rect -4301 130 -4289 1306
rect -4255 130 -4243 1306
rect -4301 118 -4243 130
rect -4123 1306 -4065 1318
rect -4123 130 -4111 1306
rect -4077 130 -4065 1306
rect -4123 118 -4065 130
rect -3945 1306 -3887 1318
rect -3945 130 -3933 1306
rect -3899 130 -3887 1306
rect -3945 118 -3887 130
rect -3767 1306 -3709 1318
rect -3767 130 -3755 1306
rect -3721 130 -3709 1306
rect -3767 118 -3709 130
rect -3589 1306 -3531 1318
rect -3589 130 -3577 1306
rect -3543 130 -3531 1306
rect -3589 118 -3531 130
rect -3411 1306 -3353 1318
rect -3411 130 -3399 1306
rect -3365 130 -3353 1306
rect -3411 118 -3353 130
rect -3233 1306 -3175 1318
rect -3233 130 -3221 1306
rect -3187 130 -3175 1306
rect -3233 118 -3175 130
rect -3055 1306 -2997 1318
rect -3055 130 -3043 1306
rect -3009 130 -2997 1306
rect -3055 118 -2997 130
rect -2877 1306 -2819 1318
rect -2877 130 -2865 1306
rect -2831 130 -2819 1306
rect -2877 118 -2819 130
rect -2699 1306 -2641 1318
rect -2699 130 -2687 1306
rect -2653 130 -2641 1306
rect -2699 118 -2641 130
rect -2521 1306 -2463 1318
rect -2521 130 -2509 1306
rect -2475 130 -2463 1306
rect -2521 118 -2463 130
rect -2343 1306 -2285 1318
rect -2343 130 -2331 1306
rect -2297 130 -2285 1306
rect -2343 118 -2285 130
rect -2165 1306 -2107 1318
rect -2165 130 -2153 1306
rect -2119 130 -2107 1306
rect -2165 118 -2107 130
rect -1987 1306 -1929 1318
rect -1987 130 -1975 1306
rect -1941 130 -1929 1306
rect -1987 118 -1929 130
rect -1809 1306 -1751 1318
rect -1809 130 -1797 1306
rect -1763 130 -1751 1306
rect -1809 118 -1751 130
rect -1631 1306 -1573 1318
rect -1631 130 -1619 1306
rect -1585 130 -1573 1306
rect -1631 118 -1573 130
rect -1453 1306 -1395 1318
rect -1453 130 -1441 1306
rect -1407 130 -1395 1306
rect -1453 118 -1395 130
rect -1275 1306 -1217 1318
rect -1275 130 -1263 1306
rect -1229 130 -1217 1306
rect -1275 118 -1217 130
rect -1097 1306 -1039 1318
rect -1097 130 -1085 1306
rect -1051 130 -1039 1306
rect -1097 118 -1039 130
rect -919 1306 -861 1318
rect -919 130 -907 1306
rect -873 130 -861 1306
rect -919 118 -861 130
rect -741 1306 -683 1318
rect -741 130 -729 1306
rect -695 130 -683 1306
rect -741 118 -683 130
rect -563 1306 -505 1318
rect -563 130 -551 1306
rect -517 130 -505 1306
rect -563 118 -505 130
rect -385 1306 -327 1318
rect -385 130 -373 1306
rect -339 130 -327 1306
rect -385 118 -327 130
rect -207 1306 -149 1318
rect -207 130 -195 1306
rect -161 130 -149 1306
rect -207 118 -149 130
rect -29 1306 29 1318
rect -29 130 -17 1306
rect 17 130 29 1306
rect -29 118 29 130
rect 149 1306 207 1318
rect 149 130 161 1306
rect 195 130 207 1306
rect 149 118 207 130
rect 327 1306 385 1318
rect 327 130 339 1306
rect 373 130 385 1306
rect 327 118 385 130
rect 505 1306 563 1318
rect 505 130 517 1306
rect 551 130 563 1306
rect 505 118 563 130
rect 683 1306 741 1318
rect 683 130 695 1306
rect 729 130 741 1306
rect 683 118 741 130
rect 861 1306 919 1318
rect 861 130 873 1306
rect 907 130 919 1306
rect 861 118 919 130
rect 1039 1306 1097 1318
rect 1039 130 1051 1306
rect 1085 130 1097 1306
rect 1039 118 1097 130
rect 1217 1306 1275 1318
rect 1217 130 1229 1306
rect 1263 130 1275 1306
rect 1217 118 1275 130
rect 1395 1306 1453 1318
rect 1395 130 1407 1306
rect 1441 130 1453 1306
rect 1395 118 1453 130
rect 1573 1306 1631 1318
rect 1573 130 1585 1306
rect 1619 130 1631 1306
rect 1573 118 1631 130
rect 1751 1306 1809 1318
rect 1751 130 1763 1306
rect 1797 130 1809 1306
rect 1751 118 1809 130
rect 1929 1306 1987 1318
rect 1929 130 1941 1306
rect 1975 130 1987 1306
rect 1929 118 1987 130
rect 2107 1306 2165 1318
rect 2107 130 2119 1306
rect 2153 130 2165 1306
rect 2107 118 2165 130
rect 2285 1306 2343 1318
rect 2285 130 2297 1306
rect 2331 130 2343 1306
rect 2285 118 2343 130
rect 2463 1306 2521 1318
rect 2463 130 2475 1306
rect 2509 130 2521 1306
rect 2463 118 2521 130
rect 2641 1306 2699 1318
rect 2641 130 2653 1306
rect 2687 130 2699 1306
rect 2641 118 2699 130
rect 2819 1306 2877 1318
rect 2819 130 2831 1306
rect 2865 130 2877 1306
rect 2819 118 2877 130
rect 2997 1306 3055 1318
rect 2997 130 3009 1306
rect 3043 130 3055 1306
rect 2997 118 3055 130
rect 3175 1306 3233 1318
rect 3175 130 3187 1306
rect 3221 130 3233 1306
rect 3175 118 3233 130
rect 3353 1306 3411 1318
rect 3353 130 3365 1306
rect 3399 130 3411 1306
rect 3353 118 3411 130
rect 3531 1306 3589 1318
rect 3531 130 3543 1306
rect 3577 130 3589 1306
rect 3531 118 3589 130
rect 3709 1306 3767 1318
rect 3709 130 3721 1306
rect 3755 130 3767 1306
rect 3709 118 3767 130
rect 3887 1306 3945 1318
rect 3887 130 3899 1306
rect 3933 130 3945 1306
rect 3887 118 3945 130
rect 4065 1306 4123 1318
rect 4065 130 4077 1306
rect 4111 130 4123 1306
rect 4065 118 4123 130
rect 4243 1306 4301 1318
rect 4243 130 4255 1306
rect 4289 130 4301 1306
rect 4243 118 4301 130
rect 4421 1306 4479 1318
rect 4421 130 4433 1306
rect 4467 130 4479 1306
rect 4421 118 4479 130
rect 4599 1306 4657 1318
rect 4599 130 4611 1306
rect 4645 130 4657 1306
rect 4599 118 4657 130
rect 4777 1306 4835 1318
rect 4777 130 4789 1306
rect 4823 130 4835 1306
rect 4777 118 4835 130
rect 4955 1306 5013 1318
rect 4955 130 4967 1306
rect 5001 130 5013 1306
rect 4955 118 5013 130
rect 5133 1306 5191 1318
rect 5133 130 5145 1306
rect 5179 130 5191 1306
rect 5133 118 5191 130
rect 5311 1306 5369 1318
rect 5311 130 5323 1306
rect 5357 130 5369 1306
rect 5311 118 5369 130
rect 5489 1306 5547 1318
rect 5489 130 5501 1306
rect 5535 130 5547 1306
rect 5489 118 5547 130
rect 5667 1306 5725 1318
rect 5667 130 5679 1306
rect 5713 130 5725 1306
rect 5667 118 5725 130
rect 5845 1306 5903 1318
rect 5845 130 5857 1306
rect 5891 130 5903 1306
rect 5845 118 5903 130
rect 6023 1306 6081 1318
rect 6023 130 6035 1306
rect 6069 130 6081 1306
rect 6023 118 6081 130
rect 6201 1306 6259 1318
rect 6201 130 6213 1306
rect 6247 130 6259 1306
rect 6201 118 6259 130
rect 6379 1306 6437 1318
rect 6379 130 6391 1306
rect 6425 130 6437 1306
rect 6379 118 6437 130
rect 6557 1306 6615 1318
rect 6557 130 6569 1306
rect 6603 130 6615 1306
rect 6557 118 6615 130
rect 6735 1306 6793 1318
rect 6735 130 6747 1306
rect 6781 130 6793 1306
rect 6735 118 6793 130
rect 6913 1306 6971 1318
rect 6913 130 6925 1306
rect 6959 130 6971 1306
rect 6913 118 6971 130
rect 7091 1306 7149 1318
rect 7091 130 7103 1306
rect 7137 130 7149 1306
rect 7091 118 7149 130
rect 7269 1306 7327 1318
rect 7269 130 7281 1306
rect 7315 130 7327 1306
rect 7269 118 7327 130
rect 7447 1306 7505 1318
rect 7447 130 7459 1306
rect 7493 130 7505 1306
rect 7447 118 7505 130
rect 7625 1306 7683 1318
rect 7625 130 7637 1306
rect 7671 130 7683 1306
rect 7625 118 7683 130
rect 7803 1306 7861 1318
rect 7803 130 7815 1306
rect 7849 130 7861 1306
rect 7803 118 7861 130
rect 7981 1306 8039 1318
rect 7981 130 7993 1306
rect 8027 130 8039 1306
rect 7981 118 8039 130
rect -8039 -130 -7981 -118
rect -8039 -1306 -8027 -130
rect -7993 -1306 -7981 -130
rect -8039 -1318 -7981 -1306
rect -7861 -130 -7803 -118
rect -7861 -1306 -7849 -130
rect -7815 -1306 -7803 -130
rect -7861 -1318 -7803 -1306
rect -7683 -130 -7625 -118
rect -7683 -1306 -7671 -130
rect -7637 -1306 -7625 -130
rect -7683 -1318 -7625 -1306
rect -7505 -130 -7447 -118
rect -7505 -1306 -7493 -130
rect -7459 -1306 -7447 -130
rect -7505 -1318 -7447 -1306
rect -7327 -130 -7269 -118
rect -7327 -1306 -7315 -130
rect -7281 -1306 -7269 -130
rect -7327 -1318 -7269 -1306
rect -7149 -130 -7091 -118
rect -7149 -1306 -7137 -130
rect -7103 -1306 -7091 -130
rect -7149 -1318 -7091 -1306
rect -6971 -130 -6913 -118
rect -6971 -1306 -6959 -130
rect -6925 -1306 -6913 -130
rect -6971 -1318 -6913 -1306
rect -6793 -130 -6735 -118
rect -6793 -1306 -6781 -130
rect -6747 -1306 -6735 -130
rect -6793 -1318 -6735 -1306
rect -6615 -130 -6557 -118
rect -6615 -1306 -6603 -130
rect -6569 -1306 -6557 -130
rect -6615 -1318 -6557 -1306
rect -6437 -130 -6379 -118
rect -6437 -1306 -6425 -130
rect -6391 -1306 -6379 -130
rect -6437 -1318 -6379 -1306
rect -6259 -130 -6201 -118
rect -6259 -1306 -6247 -130
rect -6213 -1306 -6201 -130
rect -6259 -1318 -6201 -1306
rect -6081 -130 -6023 -118
rect -6081 -1306 -6069 -130
rect -6035 -1306 -6023 -130
rect -6081 -1318 -6023 -1306
rect -5903 -130 -5845 -118
rect -5903 -1306 -5891 -130
rect -5857 -1306 -5845 -130
rect -5903 -1318 -5845 -1306
rect -5725 -130 -5667 -118
rect -5725 -1306 -5713 -130
rect -5679 -1306 -5667 -130
rect -5725 -1318 -5667 -1306
rect -5547 -130 -5489 -118
rect -5547 -1306 -5535 -130
rect -5501 -1306 -5489 -130
rect -5547 -1318 -5489 -1306
rect -5369 -130 -5311 -118
rect -5369 -1306 -5357 -130
rect -5323 -1306 -5311 -130
rect -5369 -1318 -5311 -1306
rect -5191 -130 -5133 -118
rect -5191 -1306 -5179 -130
rect -5145 -1306 -5133 -130
rect -5191 -1318 -5133 -1306
rect -5013 -130 -4955 -118
rect -5013 -1306 -5001 -130
rect -4967 -1306 -4955 -130
rect -5013 -1318 -4955 -1306
rect -4835 -130 -4777 -118
rect -4835 -1306 -4823 -130
rect -4789 -1306 -4777 -130
rect -4835 -1318 -4777 -1306
rect -4657 -130 -4599 -118
rect -4657 -1306 -4645 -130
rect -4611 -1306 -4599 -130
rect -4657 -1318 -4599 -1306
rect -4479 -130 -4421 -118
rect -4479 -1306 -4467 -130
rect -4433 -1306 -4421 -130
rect -4479 -1318 -4421 -1306
rect -4301 -130 -4243 -118
rect -4301 -1306 -4289 -130
rect -4255 -1306 -4243 -130
rect -4301 -1318 -4243 -1306
rect -4123 -130 -4065 -118
rect -4123 -1306 -4111 -130
rect -4077 -1306 -4065 -130
rect -4123 -1318 -4065 -1306
rect -3945 -130 -3887 -118
rect -3945 -1306 -3933 -130
rect -3899 -1306 -3887 -130
rect -3945 -1318 -3887 -1306
rect -3767 -130 -3709 -118
rect -3767 -1306 -3755 -130
rect -3721 -1306 -3709 -130
rect -3767 -1318 -3709 -1306
rect -3589 -130 -3531 -118
rect -3589 -1306 -3577 -130
rect -3543 -1306 -3531 -130
rect -3589 -1318 -3531 -1306
rect -3411 -130 -3353 -118
rect -3411 -1306 -3399 -130
rect -3365 -1306 -3353 -130
rect -3411 -1318 -3353 -1306
rect -3233 -130 -3175 -118
rect -3233 -1306 -3221 -130
rect -3187 -1306 -3175 -130
rect -3233 -1318 -3175 -1306
rect -3055 -130 -2997 -118
rect -3055 -1306 -3043 -130
rect -3009 -1306 -2997 -130
rect -3055 -1318 -2997 -1306
rect -2877 -130 -2819 -118
rect -2877 -1306 -2865 -130
rect -2831 -1306 -2819 -130
rect -2877 -1318 -2819 -1306
rect -2699 -130 -2641 -118
rect -2699 -1306 -2687 -130
rect -2653 -1306 -2641 -130
rect -2699 -1318 -2641 -1306
rect -2521 -130 -2463 -118
rect -2521 -1306 -2509 -130
rect -2475 -1306 -2463 -130
rect -2521 -1318 -2463 -1306
rect -2343 -130 -2285 -118
rect -2343 -1306 -2331 -130
rect -2297 -1306 -2285 -130
rect -2343 -1318 -2285 -1306
rect -2165 -130 -2107 -118
rect -2165 -1306 -2153 -130
rect -2119 -1306 -2107 -130
rect -2165 -1318 -2107 -1306
rect -1987 -130 -1929 -118
rect -1987 -1306 -1975 -130
rect -1941 -1306 -1929 -130
rect -1987 -1318 -1929 -1306
rect -1809 -130 -1751 -118
rect -1809 -1306 -1797 -130
rect -1763 -1306 -1751 -130
rect -1809 -1318 -1751 -1306
rect -1631 -130 -1573 -118
rect -1631 -1306 -1619 -130
rect -1585 -1306 -1573 -130
rect -1631 -1318 -1573 -1306
rect -1453 -130 -1395 -118
rect -1453 -1306 -1441 -130
rect -1407 -1306 -1395 -130
rect -1453 -1318 -1395 -1306
rect -1275 -130 -1217 -118
rect -1275 -1306 -1263 -130
rect -1229 -1306 -1217 -130
rect -1275 -1318 -1217 -1306
rect -1097 -130 -1039 -118
rect -1097 -1306 -1085 -130
rect -1051 -1306 -1039 -130
rect -1097 -1318 -1039 -1306
rect -919 -130 -861 -118
rect -919 -1306 -907 -130
rect -873 -1306 -861 -130
rect -919 -1318 -861 -1306
rect -741 -130 -683 -118
rect -741 -1306 -729 -130
rect -695 -1306 -683 -130
rect -741 -1318 -683 -1306
rect -563 -130 -505 -118
rect -563 -1306 -551 -130
rect -517 -1306 -505 -130
rect -563 -1318 -505 -1306
rect -385 -130 -327 -118
rect -385 -1306 -373 -130
rect -339 -1306 -327 -130
rect -385 -1318 -327 -1306
rect -207 -130 -149 -118
rect -207 -1306 -195 -130
rect -161 -1306 -149 -130
rect -207 -1318 -149 -1306
rect -29 -130 29 -118
rect -29 -1306 -17 -130
rect 17 -1306 29 -130
rect -29 -1318 29 -1306
rect 149 -130 207 -118
rect 149 -1306 161 -130
rect 195 -1306 207 -130
rect 149 -1318 207 -1306
rect 327 -130 385 -118
rect 327 -1306 339 -130
rect 373 -1306 385 -130
rect 327 -1318 385 -1306
rect 505 -130 563 -118
rect 505 -1306 517 -130
rect 551 -1306 563 -130
rect 505 -1318 563 -1306
rect 683 -130 741 -118
rect 683 -1306 695 -130
rect 729 -1306 741 -130
rect 683 -1318 741 -1306
rect 861 -130 919 -118
rect 861 -1306 873 -130
rect 907 -1306 919 -130
rect 861 -1318 919 -1306
rect 1039 -130 1097 -118
rect 1039 -1306 1051 -130
rect 1085 -1306 1097 -130
rect 1039 -1318 1097 -1306
rect 1217 -130 1275 -118
rect 1217 -1306 1229 -130
rect 1263 -1306 1275 -130
rect 1217 -1318 1275 -1306
rect 1395 -130 1453 -118
rect 1395 -1306 1407 -130
rect 1441 -1306 1453 -130
rect 1395 -1318 1453 -1306
rect 1573 -130 1631 -118
rect 1573 -1306 1585 -130
rect 1619 -1306 1631 -130
rect 1573 -1318 1631 -1306
rect 1751 -130 1809 -118
rect 1751 -1306 1763 -130
rect 1797 -1306 1809 -130
rect 1751 -1318 1809 -1306
rect 1929 -130 1987 -118
rect 1929 -1306 1941 -130
rect 1975 -1306 1987 -130
rect 1929 -1318 1987 -1306
rect 2107 -130 2165 -118
rect 2107 -1306 2119 -130
rect 2153 -1306 2165 -130
rect 2107 -1318 2165 -1306
rect 2285 -130 2343 -118
rect 2285 -1306 2297 -130
rect 2331 -1306 2343 -130
rect 2285 -1318 2343 -1306
rect 2463 -130 2521 -118
rect 2463 -1306 2475 -130
rect 2509 -1306 2521 -130
rect 2463 -1318 2521 -1306
rect 2641 -130 2699 -118
rect 2641 -1306 2653 -130
rect 2687 -1306 2699 -130
rect 2641 -1318 2699 -1306
rect 2819 -130 2877 -118
rect 2819 -1306 2831 -130
rect 2865 -1306 2877 -130
rect 2819 -1318 2877 -1306
rect 2997 -130 3055 -118
rect 2997 -1306 3009 -130
rect 3043 -1306 3055 -130
rect 2997 -1318 3055 -1306
rect 3175 -130 3233 -118
rect 3175 -1306 3187 -130
rect 3221 -1306 3233 -130
rect 3175 -1318 3233 -1306
rect 3353 -130 3411 -118
rect 3353 -1306 3365 -130
rect 3399 -1306 3411 -130
rect 3353 -1318 3411 -1306
rect 3531 -130 3589 -118
rect 3531 -1306 3543 -130
rect 3577 -1306 3589 -130
rect 3531 -1318 3589 -1306
rect 3709 -130 3767 -118
rect 3709 -1306 3721 -130
rect 3755 -1306 3767 -130
rect 3709 -1318 3767 -1306
rect 3887 -130 3945 -118
rect 3887 -1306 3899 -130
rect 3933 -1306 3945 -130
rect 3887 -1318 3945 -1306
rect 4065 -130 4123 -118
rect 4065 -1306 4077 -130
rect 4111 -1306 4123 -130
rect 4065 -1318 4123 -1306
rect 4243 -130 4301 -118
rect 4243 -1306 4255 -130
rect 4289 -1306 4301 -130
rect 4243 -1318 4301 -1306
rect 4421 -130 4479 -118
rect 4421 -1306 4433 -130
rect 4467 -1306 4479 -130
rect 4421 -1318 4479 -1306
rect 4599 -130 4657 -118
rect 4599 -1306 4611 -130
rect 4645 -1306 4657 -130
rect 4599 -1318 4657 -1306
rect 4777 -130 4835 -118
rect 4777 -1306 4789 -130
rect 4823 -1306 4835 -130
rect 4777 -1318 4835 -1306
rect 4955 -130 5013 -118
rect 4955 -1306 4967 -130
rect 5001 -1306 5013 -130
rect 4955 -1318 5013 -1306
rect 5133 -130 5191 -118
rect 5133 -1306 5145 -130
rect 5179 -1306 5191 -130
rect 5133 -1318 5191 -1306
rect 5311 -130 5369 -118
rect 5311 -1306 5323 -130
rect 5357 -1306 5369 -130
rect 5311 -1318 5369 -1306
rect 5489 -130 5547 -118
rect 5489 -1306 5501 -130
rect 5535 -1306 5547 -130
rect 5489 -1318 5547 -1306
rect 5667 -130 5725 -118
rect 5667 -1306 5679 -130
rect 5713 -1306 5725 -130
rect 5667 -1318 5725 -1306
rect 5845 -130 5903 -118
rect 5845 -1306 5857 -130
rect 5891 -1306 5903 -130
rect 5845 -1318 5903 -1306
rect 6023 -130 6081 -118
rect 6023 -1306 6035 -130
rect 6069 -1306 6081 -130
rect 6023 -1318 6081 -1306
rect 6201 -130 6259 -118
rect 6201 -1306 6213 -130
rect 6247 -1306 6259 -130
rect 6201 -1318 6259 -1306
rect 6379 -130 6437 -118
rect 6379 -1306 6391 -130
rect 6425 -1306 6437 -130
rect 6379 -1318 6437 -1306
rect 6557 -130 6615 -118
rect 6557 -1306 6569 -130
rect 6603 -1306 6615 -130
rect 6557 -1318 6615 -1306
rect 6735 -130 6793 -118
rect 6735 -1306 6747 -130
rect 6781 -1306 6793 -130
rect 6735 -1318 6793 -1306
rect 6913 -130 6971 -118
rect 6913 -1306 6925 -130
rect 6959 -1306 6971 -130
rect 6913 -1318 6971 -1306
rect 7091 -130 7149 -118
rect 7091 -1306 7103 -130
rect 7137 -1306 7149 -130
rect 7091 -1318 7149 -1306
rect 7269 -130 7327 -118
rect 7269 -1306 7281 -130
rect 7315 -1306 7327 -130
rect 7269 -1318 7327 -1306
rect 7447 -130 7505 -118
rect 7447 -1306 7459 -130
rect 7493 -1306 7505 -130
rect 7447 -1318 7505 -1306
rect 7625 -130 7683 -118
rect 7625 -1306 7637 -130
rect 7671 -1306 7683 -130
rect 7625 -1318 7683 -1306
rect 7803 -130 7861 -118
rect 7803 -1306 7815 -130
rect 7849 -1306 7861 -130
rect 7803 -1318 7861 -1306
rect 7981 -130 8039 -118
rect 7981 -1306 7993 -130
rect 8027 -1306 8039 -130
rect 7981 -1318 8039 -1306
<< pdiffc >>
rect -8027 130 -7993 1306
rect -7849 130 -7815 1306
rect -7671 130 -7637 1306
rect -7493 130 -7459 1306
rect -7315 130 -7281 1306
rect -7137 130 -7103 1306
rect -6959 130 -6925 1306
rect -6781 130 -6747 1306
rect -6603 130 -6569 1306
rect -6425 130 -6391 1306
rect -6247 130 -6213 1306
rect -6069 130 -6035 1306
rect -5891 130 -5857 1306
rect -5713 130 -5679 1306
rect -5535 130 -5501 1306
rect -5357 130 -5323 1306
rect -5179 130 -5145 1306
rect -5001 130 -4967 1306
rect -4823 130 -4789 1306
rect -4645 130 -4611 1306
rect -4467 130 -4433 1306
rect -4289 130 -4255 1306
rect -4111 130 -4077 1306
rect -3933 130 -3899 1306
rect -3755 130 -3721 1306
rect -3577 130 -3543 1306
rect -3399 130 -3365 1306
rect -3221 130 -3187 1306
rect -3043 130 -3009 1306
rect -2865 130 -2831 1306
rect -2687 130 -2653 1306
rect -2509 130 -2475 1306
rect -2331 130 -2297 1306
rect -2153 130 -2119 1306
rect -1975 130 -1941 1306
rect -1797 130 -1763 1306
rect -1619 130 -1585 1306
rect -1441 130 -1407 1306
rect -1263 130 -1229 1306
rect -1085 130 -1051 1306
rect -907 130 -873 1306
rect -729 130 -695 1306
rect -551 130 -517 1306
rect -373 130 -339 1306
rect -195 130 -161 1306
rect -17 130 17 1306
rect 161 130 195 1306
rect 339 130 373 1306
rect 517 130 551 1306
rect 695 130 729 1306
rect 873 130 907 1306
rect 1051 130 1085 1306
rect 1229 130 1263 1306
rect 1407 130 1441 1306
rect 1585 130 1619 1306
rect 1763 130 1797 1306
rect 1941 130 1975 1306
rect 2119 130 2153 1306
rect 2297 130 2331 1306
rect 2475 130 2509 1306
rect 2653 130 2687 1306
rect 2831 130 2865 1306
rect 3009 130 3043 1306
rect 3187 130 3221 1306
rect 3365 130 3399 1306
rect 3543 130 3577 1306
rect 3721 130 3755 1306
rect 3899 130 3933 1306
rect 4077 130 4111 1306
rect 4255 130 4289 1306
rect 4433 130 4467 1306
rect 4611 130 4645 1306
rect 4789 130 4823 1306
rect 4967 130 5001 1306
rect 5145 130 5179 1306
rect 5323 130 5357 1306
rect 5501 130 5535 1306
rect 5679 130 5713 1306
rect 5857 130 5891 1306
rect 6035 130 6069 1306
rect 6213 130 6247 1306
rect 6391 130 6425 1306
rect 6569 130 6603 1306
rect 6747 130 6781 1306
rect 6925 130 6959 1306
rect 7103 130 7137 1306
rect 7281 130 7315 1306
rect 7459 130 7493 1306
rect 7637 130 7671 1306
rect 7815 130 7849 1306
rect 7993 130 8027 1306
rect -8027 -1306 -7993 -130
rect -7849 -1306 -7815 -130
rect -7671 -1306 -7637 -130
rect -7493 -1306 -7459 -130
rect -7315 -1306 -7281 -130
rect -7137 -1306 -7103 -130
rect -6959 -1306 -6925 -130
rect -6781 -1306 -6747 -130
rect -6603 -1306 -6569 -130
rect -6425 -1306 -6391 -130
rect -6247 -1306 -6213 -130
rect -6069 -1306 -6035 -130
rect -5891 -1306 -5857 -130
rect -5713 -1306 -5679 -130
rect -5535 -1306 -5501 -130
rect -5357 -1306 -5323 -130
rect -5179 -1306 -5145 -130
rect -5001 -1306 -4967 -130
rect -4823 -1306 -4789 -130
rect -4645 -1306 -4611 -130
rect -4467 -1306 -4433 -130
rect -4289 -1306 -4255 -130
rect -4111 -1306 -4077 -130
rect -3933 -1306 -3899 -130
rect -3755 -1306 -3721 -130
rect -3577 -1306 -3543 -130
rect -3399 -1306 -3365 -130
rect -3221 -1306 -3187 -130
rect -3043 -1306 -3009 -130
rect -2865 -1306 -2831 -130
rect -2687 -1306 -2653 -130
rect -2509 -1306 -2475 -130
rect -2331 -1306 -2297 -130
rect -2153 -1306 -2119 -130
rect -1975 -1306 -1941 -130
rect -1797 -1306 -1763 -130
rect -1619 -1306 -1585 -130
rect -1441 -1306 -1407 -130
rect -1263 -1306 -1229 -130
rect -1085 -1306 -1051 -130
rect -907 -1306 -873 -130
rect -729 -1306 -695 -130
rect -551 -1306 -517 -130
rect -373 -1306 -339 -130
rect -195 -1306 -161 -130
rect -17 -1306 17 -130
rect 161 -1306 195 -130
rect 339 -1306 373 -130
rect 517 -1306 551 -130
rect 695 -1306 729 -130
rect 873 -1306 907 -130
rect 1051 -1306 1085 -130
rect 1229 -1306 1263 -130
rect 1407 -1306 1441 -130
rect 1585 -1306 1619 -130
rect 1763 -1306 1797 -130
rect 1941 -1306 1975 -130
rect 2119 -1306 2153 -130
rect 2297 -1306 2331 -130
rect 2475 -1306 2509 -130
rect 2653 -1306 2687 -130
rect 2831 -1306 2865 -130
rect 3009 -1306 3043 -130
rect 3187 -1306 3221 -130
rect 3365 -1306 3399 -130
rect 3543 -1306 3577 -130
rect 3721 -1306 3755 -130
rect 3899 -1306 3933 -130
rect 4077 -1306 4111 -130
rect 4255 -1306 4289 -130
rect 4433 -1306 4467 -130
rect 4611 -1306 4645 -130
rect 4789 -1306 4823 -130
rect 4967 -1306 5001 -130
rect 5145 -1306 5179 -130
rect 5323 -1306 5357 -130
rect 5501 -1306 5535 -130
rect 5679 -1306 5713 -130
rect 5857 -1306 5891 -130
rect 6035 -1306 6069 -130
rect 6213 -1306 6247 -130
rect 6391 -1306 6425 -130
rect 6569 -1306 6603 -130
rect 6747 -1306 6781 -130
rect 6925 -1306 6959 -130
rect 7103 -1306 7137 -130
rect 7281 -1306 7315 -130
rect 7459 -1306 7493 -130
rect 7637 -1306 7671 -130
rect 7815 -1306 7849 -130
rect 7993 -1306 8027 -130
<< nsubdiff >>
rect -8141 1467 -8045 1501
rect 8045 1467 8141 1501
rect -8141 1405 -8107 1467
rect 8107 1405 8141 1467
rect -8141 -1467 -8107 -1405
rect 8107 -1467 8141 -1405
rect -8141 -1501 -8045 -1467
rect 8045 -1501 8141 -1467
<< nsubdiffcont >>
rect -8045 1467 8045 1501
rect -8141 -1405 -8107 1405
rect 8107 -1405 8141 1405
rect -8045 -1501 8045 -1467
<< poly >>
rect -7981 1399 -7861 1415
rect -7981 1365 -7965 1399
rect -7877 1365 -7861 1399
rect -7981 1318 -7861 1365
rect -7803 1399 -7683 1415
rect -7803 1365 -7787 1399
rect -7699 1365 -7683 1399
rect -7803 1318 -7683 1365
rect -7625 1399 -7505 1415
rect -7625 1365 -7609 1399
rect -7521 1365 -7505 1399
rect -7625 1318 -7505 1365
rect -7447 1399 -7327 1415
rect -7447 1365 -7431 1399
rect -7343 1365 -7327 1399
rect -7447 1318 -7327 1365
rect -7269 1399 -7149 1415
rect -7269 1365 -7253 1399
rect -7165 1365 -7149 1399
rect -7269 1318 -7149 1365
rect -7091 1399 -6971 1415
rect -7091 1365 -7075 1399
rect -6987 1365 -6971 1399
rect -7091 1318 -6971 1365
rect -6913 1399 -6793 1415
rect -6913 1365 -6897 1399
rect -6809 1365 -6793 1399
rect -6913 1318 -6793 1365
rect -6735 1399 -6615 1415
rect -6735 1365 -6719 1399
rect -6631 1365 -6615 1399
rect -6735 1318 -6615 1365
rect -6557 1399 -6437 1415
rect -6557 1365 -6541 1399
rect -6453 1365 -6437 1399
rect -6557 1318 -6437 1365
rect -6379 1399 -6259 1415
rect -6379 1365 -6363 1399
rect -6275 1365 -6259 1399
rect -6379 1318 -6259 1365
rect -6201 1399 -6081 1415
rect -6201 1365 -6185 1399
rect -6097 1365 -6081 1399
rect -6201 1318 -6081 1365
rect -6023 1399 -5903 1415
rect -6023 1365 -6007 1399
rect -5919 1365 -5903 1399
rect -6023 1318 -5903 1365
rect -5845 1399 -5725 1415
rect -5845 1365 -5829 1399
rect -5741 1365 -5725 1399
rect -5845 1318 -5725 1365
rect -5667 1399 -5547 1415
rect -5667 1365 -5651 1399
rect -5563 1365 -5547 1399
rect -5667 1318 -5547 1365
rect -5489 1399 -5369 1415
rect -5489 1365 -5473 1399
rect -5385 1365 -5369 1399
rect -5489 1318 -5369 1365
rect -5311 1399 -5191 1415
rect -5311 1365 -5295 1399
rect -5207 1365 -5191 1399
rect -5311 1318 -5191 1365
rect -5133 1399 -5013 1415
rect -5133 1365 -5117 1399
rect -5029 1365 -5013 1399
rect -5133 1318 -5013 1365
rect -4955 1399 -4835 1415
rect -4955 1365 -4939 1399
rect -4851 1365 -4835 1399
rect -4955 1318 -4835 1365
rect -4777 1399 -4657 1415
rect -4777 1365 -4761 1399
rect -4673 1365 -4657 1399
rect -4777 1318 -4657 1365
rect -4599 1399 -4479 1415
rect -4599 1365 -4583 1399
rect -4495 1365 -4479 1399
rect -4599 1318 -4479 1365
rect -4421 1399 -4301 1415
rect -4421 1365 -4405 1399
rect -4317 1365 -4301 1399
rect -4421 1318 -4301 1365
rect -4243 1399 -4123 1415
rect -4243 1365 -4227 1399
rect -4139 1365 -4123 1399
rect -4243 1318 -4123 1365
rect -4065 1399 -3945 1415
rect -4065 1365 -4049 1399
rect -3961 1365 -3945 1399
rect -4065 1318 -3945 1365
rect -3887 1399 -3767 1415
rect -3887 1365 -3871 1399
rect -3783 1365 -3767 1399
rect -3887 1318 -3767 1365
rect -3709 1399 -3589 1415
rect -3709 1365 -3693 1399
rect -3605 1365 -3589 1399
rect -3709 1318 -3589 1365
rect -3531 1399 -3411 1415
rect -3531 1365 -3515 1399
rect -3427 1365 -3411 1399
rect -3531 1318 -3411 1365
rect -3353 1399 -3233 1415
rect -3353 1365 -3337 1399
rect -3249 1365 -3233 1399
rect -3353 1318 -3233 1365
rect -3175 1399 -3055 1415
rect -3175 1365 -3159 1399
rect -3071 1365 -3055 1399
rect -3175 1318 -3055 1365
rect -2997 1399 -2877 1415
rect -2997 1365 -2981 1399
rect -2893 1365 -2877 1399
rect -2997 1318 -2877 1365
rect -2819 1399 -2699 1415
rect -2819 1365 -2803 1399
rect -2715 1365 -2699 1399
rect -2819 1318 -2699 1365
rect -2641 1399 -2521 1415
rect -2641 1365 -2625 1399
rect -2537 1365 -2521 1399
rect -2641 1318 -2521 1365
rect -2463 1399 -2343 1415
rect -2463 1365 -2447 1399
rect -2359 1365 -2343 1399
rect -2463 1318 -2343 1365
rect -2285 1399 -2165 1415
rect -2285 1365 -2269 1399
rect -2181 1365 -2165 1399
rect -2285 1318 -2165 1365
rect -2107 1399 -1987 1415
rect -2107 1365 -2091 1399
rect -2003 1365 -1987 1399
rect -2107 1318 -1987 1365
rect -1929 1399 -1809 1415
rect -1929 1365 -1913 1399
rect -1825 1365 -1809 1399
rect -1929 1318 -1809 1365
rect -1751 1399 -1631 1415
rect -1751 1365 -1735 1399
rect -1647 1365 -1631 1399
rect -1751 1318 -1631 1365
rect -1573 1399 -1453 1415
rect -1573 1365 -1557 1399
rect -1469 1365 -1453 1399
rect -1573 1318 -1453 1365
rect -1395 1399 -1275 1415
rect -1395 1365 -1379 1399
rect -1291 1365 -1275 1399
rect -1395 1318 -1275 1365
rect -1217 1399 -1097 1415
rect -1217 1365 -1201 1399
rect -1113 1365 -1097 1399
rect -1217 1318 -1097 1365
rect -1039 1399 -919 1415
rect -1039 1365 -1023 1399
rect -935 1365 -919 1399
rect -1039 1318 -919 1365
rect -861 1399 -741 1415
rect -861 1365 -845 1399
rect -757 1365 -741 1399
rect -861 1318 -741 1365
rect -683 1399 -563 1415
rect -683 1365 -667 1399
rect -579 1365 -563 1399
rect -683 1318 -563 1365
rect -505 1399 -385 1415
rect -505 1365 -489 1399
rect -401 1365 -385 1399
rect -505 1318 -385 1365
rect -327 1399 -207 1415
rect -327 1365 -311 1399
rect -223 1365 -207 1399
rect -327 1318 -207 1365
rect -149 1399 -29 1415
rect -149 1365 -133 1399
rect -45 1365 -29 1399
rect -149 1318 -29 1365
rect 29 1399 149 1415
rect 29 1365 45 1399
rect 133 1365 149 1399
rect 29 1318 149 1365
rect 207 1399 327 1415
rect 207 1365 223 1399
rect 311 1365 327 1399
rect 207 1318 327 1365
rect 385 1399 505 1415
rect 385 1365 401 1399
rect 489 1365 505 1399
rect 385 1318 505 1365
rect 563 1399 683 1415
rect 563 1365 579 1399
rect 667 1365 683 1399
rect 563 1318 683 1365
rect 741 1399 861 1415
rect 741 1365 757 1399
rect 845 1365 861 1399
rect 741 1318 861 1365
rect 919 1399 1039 1415
rect 919 1365 935 1399
rect 1023 1365 1039 1399
rect 919 1318 1039 1365
rect 1097 1399 1217 1415
rect 1097 1365 1113 1399
rect 1201 1365 1217 1399
rect 1097 1318 1217 1365
rect 1275 1399 1395 1415
rect 1275 1365 1291 1399
rect 1379 1365 1395 1399
rect 1275 1318 1395 1365
rect 1453 1399 1573 1415
rect 1453 1365 1469 1399
rect 1557 1365 1573 1399
rect 1453 1318 1573 1365
rect 1631 1399 1751 1415
rect 1631 1365 1647 1399
rect 1735 1365 1751 1399
rect 1631 1318 1751 1365
rect 1809 1399 1929 1415
rect 1809 1365 1825 1399
rect 1913 1365 1929 1399
rect 1809 1318 1929 1365
rect 1987 1399 2107 1415
rect 1987 1365 2003 1399
rect 2091 1365 2107 1399
rect 1987 1318 2107 1365
rect 2165 1399 2285 1415
rect 2165 1365 2181 1399
rect 2269 1365 2285 1399
rect 2165 1318 2285 1365
rect 2343 1399 2463 1415
rect 2343 1365 2359 1399
rect 2447 1365 2463 1399
rect 2343 1318 2463 1365
rect 2521 1399 2641 1415
rect 2521 1365 2537 1399
rect 2625 1365 2641 1399
rect 2521 1318 2641 1365
rect 2699 1399 2819 1415
rect 2699 1365 2715 1399
rect 2803 1365 2819 1399
rect 2699 1318 2819 1365
rect 2877 1399 2997 1415
rect 2877 1365 2893 1399
rect 2981 1365 2997 1399
rect 2877 1318 2997 1365
rect 3055 1399 3175 1415
rect 3055 1365 3071 1399
rect 3159 1365 3175 1399
rect 3055 1318 3175 1365
rect 3233 1399 3353 1415
rect 3233 1365 3249 1399
rect 3337 1365 3353 1399
rect 3233 1318 3353 1365
rect 3411 1399 3531 1415
rect 3411 1365 3427 1399
rect 3515 1365 3531 1399
rect 3411 1318 3531 1365
rect 3589 1399 3709 1415
rect 3589 1365 3605 1399
rect 3693 1365 3709 1399
rect 3589 1318 3709 1365
rect 3767 1399 3887 1415
rect 3767 1365 3783 1399
rect 3871 1365 3887 1399
rect 3767 1318 3887 1365
rect 3945 1399 4065 1415
rect 3945 1365 3961 1399
rect 4049 1365 4065 1399
rect 3945 1318 4065 1365
rect 4123 1399 4243 1415
rect 4123 1365 4139 1399
rect 4227 1365 4243 1399
rect 4123 1318 4243 1365
rect 4301 1399 4421 1415
rect 4301 1365 4317 1399
rect 4405 1365 4421 1399
rect 4301 1318 4421 1365
rect 4479 1399 4599 1415
rect 4479 1365 4495 1399
rect 4583 1365 4599 1399
rect 4479 1318 4599 1365
rect 4657 1399 4777 1415
rect 4657 1365 4673 1399
rect 4761 1365 4777 1399
rect 4657 1318 4777 1365
rect 4835 1399 4955 1415
rect 4835 1365 4851 1399
rect 4939 1365 4955 1399
rect 4835 1318 4955 1365
rect 5013 1399 5133 1415
rect 5013 1365 5029 1399
rect 5117 1365 5133 1399
rect 5013 1318 5133 1365
rect 5191 1399 5311 1415
rect 5191 1365 5207 1399
rect 5295 1365 5311 1399
rect 5191 1318 5311 1365
rect 5369 1399 5489 1415
rect 5369 1365 5385 1399
rect 5473 1365 5489 1399
rect 5369 1318 5489 1365
rect 5547 1399 5667 1415
rect 5547 1365 5563 1399
rect 5651 1365 5667 1399
rect 5547 1318 5667 1365
rect 5725 1399 5845 1415
rect 5725 1365 5741 1399
rect 5829 1365 5845 1399
rect 5725 1318 5845 1365
rect 5903 1399 6023 1415
rect 5903 1365 5919 1399
rect 6007 1365 6023 1399
rect 5903 1318 6023 1365
rect 6081 1399 6201 1415
rect 6081 1365 6097 1399
rect 6185 1365 6201 1399
rect 6081 1318 6201 1365
rect 6259 1399 6379 1415
rect 6259 1365 6275 1399
rect 6363 1365 6379 1399
rect 6259 1318 6379 1365
rect 6437 1399 6557 1415
rect 6437 1365 6453 1399
rect 6541 1365 6557 1399
rect 6437 1318 6557 1365
rect 6615 1399 6735 1415
rect 6615 1365 6631 1399
rect 6719 1365 6735 1399
rect 6615 1318 6735 1365
rect 6793 1399 6913 1415
rect 6793 1365 6809 1399
rect 6897 1365 6913 1399
rect 6793 1318 6913 1365
rect 6971 1399 7091 1415
rect 6971 1365 6987 1399
rect 7075 1365 7091 1399
rect 6971 1318 7091 1365
rect 7149 1399 7269 1415
rect 7149 1365 7165 1399
rect 7253 1365 7269 1399
rect 7149 1318 7269 1365
rect 7327 1399 7447 1415
rect 7327 1365 7343 1399
rect 7431 1365 7447 1399
rect 7327 1318 7447 1365
rect 7505 1399 7625 1415
rect 7505 1365 7521 1399
rect 7609 1365 7625 1399
rect 7505 1318 7625 1365
rect 7683 1399 7803 1415
rect 7683 1365 7699 1399
rect 7787 1365 7803 1399
rect 7683 1318 7803 1365
rect 7861 1399 7981 1415
rect 7861 1365 7877 1399
rect 7965 1365 7981 1399
rect 7861 1318 7981 1365
rect -7981 71 -7861 118
rect -7981 37 -7965 71
rect -7877 37 -7861 71
rect -7981 21 -7861 37
rect -7803 71 -7683 118
rect -7803 37 -7787 71
rect -7699 37 -7683 71
rect -7803 21 -7683 37
rect -7625 71 -7505 118
rect -7625 37 -7609 71
rect -7521 37 -7505 71
rect -7625 21 -7505 37
rect -7447 71 -7327 118
rect -7447 37 -7431 71
rect -7343 37 -7327 71
rect -7447 21 -7327 37
rect -7269 71 -7149 118
rect -7269 37 -7253 71
rect -7165 37 -7149 71
rect -7269 21 -7149 37
rect -7091 71 -6971 118
rect -7091 37 -7075 71
rect -6987 37 -6971 71
rect -7091 21 -6971 37
rect -6913 71 -6793 118
rect -6913 37 -6897 71
rect -6809 37 -6793 71
rect -6913 21 -6793 37
rect -6735 71 -6615 118
rect -6735 37 -6719 71
rect -6631 37 -6615 71
rect -6735 21 -6615 37
rect -6557 71 -6437 118
rect -6557 37 -6541 71
rect -6453 37 -6437 71
rect -6557 21 -6437 37
rect -6379 71 -6259 118
rect -6379 37 -6363 71
rect -6275 37 -6259 71
rect -6379 21 -6259 37
rect -6201 71 -6081 118
rect -6201 37 -6185 71
rect -6097 37 -6081 71
rect -6201 21 -6081 37
rect -6023 71 -5903 118
rect -6023 37 -6007 71
rect -5919 37 -5903 71
rect -6023 21 -5903 37
rect -5845 71 -5725 118
rect -5845 37 -5829 71
rect -5741 37 -5725 71
rect -5845 21 -5725 37
rect -5667 71 -5547 118
rect -5667 37 -5651 71
rect -5563 37 -5547 71
rect -5667 21 -5547 37
rect -5489 71 -5369 118
rect -5489 37 -5473 71
rect -5385 37 -5369 71
rect -5489 21 -5369 37
rect -5311 71 -5191 118
rect -5311 37 -5295 71
rect -5207 37 -5191 71
rect -5311 21 -5191 37
rect -5133 71 -5013 118
rect -5133 37 -5117 71
rect -5029 37 -5013 71
rect -5133 21 -5013 37
rect -4955 71 -4835 118
rect -4955 37 -4939 71
rect -4851 37 -4835 71
rect -4955 21 -4835 37
rect -4777 71 -4657 118
rect -4777 37 -4761 71
rect -4673 37 -4657 71
rect -4777 21 -4657 37
rect -4599 71 -4479 118
rect -4599 37 -4583 71
rect -4495 37 -4479 71
rect -4599 21 -4479 37
rect -4421 71 -4301 118
rect -4421 37 -4405 71
rect -4317 37 -4301 71
rect -4421 21 -4301 37
rect -4243 71 -4123 118
rect -4243 37 -4227 71
rect -4139 37 -4123 71
rect -4243 21 -4123 37
rect -4065 71 -3945 118
rect -4065 37 -4049 71
rect -3961 37 -3945 71
rect -4065 21 -3945 37
rect -3887 71 -3767 118
rect -3887 37 -3871 71
rect -3783 37 -3767 71
rect -3887 21 -3767 37
rect -3709 71 -3589 118
rect -3709 37 -3693 71
rect -3605 37 -3589 71
rect -3709 21 -3589 37
rect -3531 71 -3411 118
rect -3531 37 -3515 71
rect -3427 37 -3411 71
rect -3531 21 -3411 37
rect -3353 71 -3233 118
rect -3353 37 -3337 71
rect -3249 37 -3233 71
rect -3353 21 -3233 37
rect -3175 71 -3055 118
rect -3175 37 -3159 71
rect -3071 37 -3055 71
rect -3175 21 -3055 37
rect -2997 71 -2877 118
rect -2997 37 -2981 71
rect -2893 37 -2877 71
rect -2997 21 -2877 37
rect -2819 71 -2699 118
rect -2819 37 -2803 71
rect -2715 37 -2699 71
rect -2819 21 -2699 37
rect -2641 71 -2521 118
rect -2641 37 -2625 71
rect -2537 37 -2521 71
rect -2641 21 -2521 37
rect -2463 71 -2343 118
rect -2463 37 -2447 71
rect -2359 37 -2343 71
rect -2463 21 -2343 37
rect -2285 71 -2165 118
rect -2285 37 -2269 71
rect -2181 37 -2165 71
rect -2285 21 -2165 37
rect -2107 71 -1987 118
rect -2107 37 -2091 71
rect -2003 37 -1987 71
rect -2107 21 -1987 37
rect -1929 71 -1809 118
rect -1929 37 -1913 71
rect -1825 37 -1809 71
rect -1929 21 -1809 37
rect -1751 71 -1631 118
rect -1751 37 -1735 71
rect -1647 37 -1631 71
rect -1751 21 -1631 37
rect -1573 71 -1453 118
rect -1573 37 -1557 71
rect -1469 37 -1453 71
rect -1573 21 -1453 37
rect -1395 71 -1275 118
rect -1395 37 -1379 71
rect -1291 37 -1275 71
rect -1395 21 -1275 37
rect -1217 71 -1097 118
rect -1217 37 -1201 71
rect -1113 37 -1097 71
rect -1217 21 -1097 37
rect -1039 71 -919 118
rect -1039 37 -1023 71
rect -935 37 -919 71
rect -1039 21 -919 37
rect -861 71 -741 118
rect -861 37 -845 71
rect -757 37 -741 71
rect -861 21 -741 37
rect -683 71 -563 118
rect -683 37 -667 71
rect -579 37 -563 71
rect -683 21 -563 37
rect -505 71 -385 118
rect -505 37 -489 71
rect -401 37 -385 71
rect -505 21 -385 37
rect -327 71 -207 118
rect -327 37 -311 71
rect -223 37 -207 71
rect -327 21 -207 37
rect -149 71 -29 118
rect -149 37 -133 71
rect -45 37 -29 71
rect -149 21 -29 37
rect 29 71 149 118
rect 29 37 45 71
rect 133 37 149 71
rect 29 21 149 37
rect 207 71 327 118
rect 207 37 223 71
rect 311 37 327 71
rect 207 21 327 37
rect 385 71 505 118
rect 385 37 401 71
rect 489 37 505 71
rect 385 21 505 37
rect 563 71 683 118
rect 563 37 579 71
rect 667 37 683 71
rect 563 21 683 37
rect 741 71 861 118
rect 741 37 757 71
rect 845 37 861 71
rect 741 21 861 37
rect 919 71 1039 118
rect 919 37 935 71
rect 1023 37 1039 71
rect 919 21 1039 37
rect 1097 71 1217 118
rect 1097 37 1113 71
rect 1201 37 1217 71
rect 1097 21 1217 37
rect 1275 71 1395 118
rect 1275 37 1291 71
rect 1379 37 1395 71
rect 1275 21 1395 37
rect 1453 71 1573 118
rect 1453 37 1469 71
rect 1557 37 1573 71
rect 1453 21 1573 37
rect 1631 71 1751 118
rect 1631 37 1647 71
rect 1735 37 1751 71
rect 1631 21 1751 37
rect 1809 71 1929 118
rect 1809 37 1825 71
rect 1913 37 1929 71
rect 1809 21 1929 37
rect 1987 71 2107 118
rect 1987 37 2003 71
rect 2091 37 2107 71
rect 1987 21 2107 37
rect 2165 71 2285 118
rect 2165 37 2181 71
rect 2269 37 2285 71
rect 2165 21 2285 37
rect 2343 71 2463 118
rect 2343 37 2359 71
rect 2447 37 2463 71
rect 2343 21 2463 37
rect 2521 71 2641 118
rect 2521 37 2537 71
rect 2625 37 2641 71
rect 2521 21 2641 37
rect 2699 71 2819 118
rect 2699 37 2715 71
rect 2803 37 2819 71
rect 2699 21 2819 37
rect 2877 71 2997 118
rect 2877 37 2893 71
rect 2981 37 2997 71
rect 2877 21 2997 37
rect 3055 71 3175 118
rect 3055 37 3071 71
rect 3159 37 3175 71
rect 3055 21 3175 37
rect 3233 71 3353 118
rect 3233 37 3249 71
rect 3337 37 3353 71
rect 3233 21 3353 37
rect 3411 71 3531 118
rect 3411 37 3427 71
rect 3515 37 3531 71
rect 3411 21 3531 37
rect 3589 71 3709 118
rect 3589 37 3605 71
rect 3693 37 3709 71
rect 3589 21 3709 37
rect 3767 71 3887 118
rect 3767 37 3783 71
rect 3871 37 3887 71
rect 3767 21 3887 37
rect 3945 71 4065 118
rect 3945 37 3961 71
rect 4049 37 4065 71
rect 3945 21 4065 37
rect 4123 71 4243 118
rect 4123 37 4139 71
rect 4227 37 4243 71
rect 4123 21 4243 37
rect 4301 71 4421 118
rect 4301 37 4317 71
rect 4405 37 4421 71
rect 4301 21 4421 37
rect 4479 71 4599 118
rect 4479 37 4495 71
rect 4583 37 4599 71
rect 4479 21 4599 37
rect 4657 71 4777 118
rect 4657 37 4673 71
rect 4761 37 4777 71
rect 4657 21 4777 37
rect 4835 71 4955 118
rect 4835 37 4851 71
rect 4939 37 4955 71
rect 4835 21 4955 37
rect 5013 71 5133 118
rect 5013 37 5029 71
rect 5117 37 5133 71
rect 5013 21 5133 37
rect 5191 71 5311 118
rect 5191 37 5207 71
rect 5295 37 5311 71
rect 5191 21 5311 37
rect 5369 71 5489 118
rect 5369 37 5385 71
rect 5473 37 5489 71
rect 5369 21 5489 37
rect 5547 71 5667 118
rect 5547 37 5563 71
rect 5651 37 5667 71
rect 5547 21 5667 37
rect 5725 71 5845 118
rect 5725 37 5741 71
rect 5829 37 5845 71
rect 5725 21 5845 37
rect 5903 71 6023 118
rect 5903 37 5919 71
rect 6007 37 6023 71
rect 5903 21 6023 37
rect 6081 71 6201 118
rect 6081 37 6097 71
rect 6185 37 6201 71
rect 6081 21 6201 37
rect 6259 71 6379 118
rect 6259 37 6275 71
rect 6363 37 6379 71
rect 6259 21 6379 37
rect 6437 71 6557 118
rect 6437 37 6453 71
rect 6541 37 6557 71
rect 6437 21 6557 37
rect 6615 71 6735 118
rect 6615 37 6631 71
rect 6719 37 6735 71
rect 6615 21 6735 37
rect 6793 71 6913 118
rect 6793 37 6809 71
rect 6897 37 6913 71
rect 6793 21 6913 37
rect 6971 71 7091 118
rect 6971 37 6987 71
rect 7075 37 7091 71
rect 6971 21 7091 37
rect 7149 71 7269 118
rect 7149 37 7165 71
rect 7253 37 7269 71
rect 7149 21 7269 37
rect 7327 71 7447 118
rect 7327 37 7343 71
rect 7431 37 7447 71
rect 7327 21 7447 37
rect 7505 71 7625 118
rect 7505 37 7521 71
rect 7609 37 7625 71
rect 7505 21 7625 37
rect 7683 71 7803 118
rect 7683 37 7699 71
rect 7787 37 7803 71
rect 7683 21 7803 37
rect 7861 71 7981 118
rect 7861 37 7877 71
rect 7965 37 7981 71
rect 7861 21 7981 37
rect -7981 -37 -7861 -21
rect -7981 -71 -7965 -37
rect -7877 -71 -7861 -37
rect -7981 -118 -7861 -71
rect -7803 -37 -7683 -21
rect -7803 -71 -7787 -37
rect -7699 -71 -7683 -37
rect -7803 -118 -7683 -71
rect -7625 -37 -7505 -21
rect -7625 -71 -7609 -37
rect -7521 -71 -7505 -37
rect -7625 -118 -7505 -71
rect -7447 -37 -7327 -21
rect -7447 -71 -7431 -37
rect -7343 -71 -7327 -37
rect -7447 -118 -7327 -71
rect -7269 -37 -7149 -21
rect -7269 -71 -7253 -37
rect -7165 -71 -7149 -37
rect -7269 -118 -7149 -71
rect -7091 -37 -6971 -21
rect -7091 -71 -7075 -37
rect -6987 -71 -6971 -37
rect -7091 -118 -6971 -71
rect -6913 -37 -6793 -21
rect -6913 -71 -6897 -37
rect -6809 -71 -6793 -37
rect -6913 -118 -6793 -71
rect -6735 -37 -6615 -21
rect -6735 -71 -6719 -37
rect -6631 -71 -6615 -37
rect -6735 -118 -6615 -71
rect -6557 -37 -6437 -21
rect -6557 -71 -6541 -37
rect -6453 -71 -6437 -37
rect -6557 -118 -6437 -71
rect -6379 -37 -6259 -21
rect -6379 -71 -6363 -37
rect -6275 -71 -6259 -37
rect -6379 -118 -6259 -71
rect -6201 -37 -6081 -21
rect -6201 -71 -6185 -37
rect -6097 -71 -6081 -37
rect -6201 -118 -6081 -71
rect -6023 -37 -5903 -21
rect -6023 -71 -6007 -37
rect -5919 -71 -5903 -37
rect -6023 -118 -5903 -71
rect -5845 -37 -5725 -21
rect -5845 -71 -5829 -37
rect -5741 -71 -5725 -37
rect -5845 -118 -5725 -71
rect -5667 -37 -5547 -21
rect -5667 -71 -5651 -37
rect -5563 -71 -5547 -37
rect -5667 -118 -5547 -71
rect -5489 -37 -5369 -21
rect -5489 -71 -5473 -37
rect -5385 -71 -5369 -37
rect -5489 -118 -5369 -71
rect -5311 -37 -5191 -21
rect -5311 -71 -5295 -37
rect -5207 -71 -5191 -37
rect -5311 -118 -5191 -71
rect -5133 -37 -5013 -21
rect -5133 -71 -5117 -37
rect -5029 -71 -5013 -37
rect -5133 -118 -5013 -71
rect -4955 -37 -4835 -21
rect -4955 -71 -4939 -37
rect -4851 -71 -4835 -37
rect -4955 -118 -4835 -71
rect -4777 -37 -4657 -21
rect -4777 -71 -4761 -37
rect -4673 -71 -4657 -37
rect -4777 -118 -4657 -71
rect -4599 -37 -4479 -21
rect -4599 -71 -4583 -37
rect -4495 -71 -4479 -37
rect -4599 -118 -4479 -71
rect -4421 -37 -4301 -21
rect -4421 -71 -4405 -37
rect -4317 -71 -4301 -37
rect -4421 -118 -4301 -71
rect -4243 -37 -4123 -21
rect -4243 -71 -4227 -37
rect -4139 -71 -4123 -37
rect -4243 -118 -4123 -71
rect -4065 -37 -3945 -21
rect -4065 -71 -4049 -37
rect -3961 -71 -3945 -37
rect -4065 -118 -3945 -71
rect -3887 -37 -3767 -21
rect -3887 -71 -3871 -37
rect -3783 -71 -3767 -37
rect -3887 -118 -3767 -71
rect -3709 -37 -3589 -21
rect -3709 -71 -3693 -37
rect -3605 -71 -3589 -37
rect -3709 -118 -3589 -71
rect -3531 -37 -3411 -21
rect -3531 -71 -3515 -37
rect -3427 -71 -3411 -37
rect -3531 -118 -3411 -71
rect -3353 -37 -3233 -21
rect -3353 -71 -3337 -37
rect -3249 -71 -3233 -37
rect -3353 -118 -3233 -71
rect -3175 -37 -3055 -21
rect -3175 -71 -3159 -37
rect -3071 -71 -3055 -37
rect -3175 -118 -3055 -71
rect -2997 -37 -2877 -21
rect -2997 -71 -2981 -37
rect -2893 -71 -2877 -37
rect -2997 -118 -2877 -71
rect -2819 -37 -2699 -21
rect -2819 -71 -2803 -37
rect -2715 -71 -2699 -37
rect -2819 -118 -2699 -71
rect -2641 -37 -2521 -21
rect -2641 -71 -2625 -37
rect -2537 -71 -2521 -37
rect -2641 -118 -2521 -71
rect -2463 -37 -2343 -21
rect -2463 -71 -2447 -37
rect -2359 -71 -2343 -37
rect -2463 -118 -2343 -71
rect -2285 -37 -2165 -21
rect -2285 -71 -2269 -37
rect -2181 -71 -2165 -37
rect -2285 -118 -2165 -71
rect -2107 -37 -1987 -21
rect -2107 -71 -2091 -37
rect -2003 -71 -1987 -37
rect -2107 -118 -1987 -71
rect -1929 -37 -1809 -21
rect -1929 -71 -1913 -37
rect -1825 -71 -1809 -37
rect -1929 -118 -1809 -71
rect -1751 -37 -1631 -21
rect -1751 -71 -1735 -37
rect -1647 -71 -1631 -37
rect -1751 -118 -1631 -71
rect -1573 -37 -1453 -21
rect -1573 -71 -1557 -37
rect -1469 -71 -1453 -37
rect -1573 -118 -1453 -71
rect -1395 -37 -1275 -21
rect -1395 -71 -1379 -37
rect -1291 -71 -1275 -37
rect -1395 -118 -1275 -71
rect -1217 -37 -1097 -21
rect -1217 -71 -1201 -37
rect -1113 -71 -1097 -37
rect -1217 -118 -1097 -71
rect -1039 -37 -919 -21
rect -1039 -71 -1023 -37
rect -935 -71 -919 -37
rect -1039 -118 -919 -71
rect -861 -37 -741 -21
rect -861 -71 -845 -37
rect -757 -71 -741 -37
rect -861 -118 -741 -71
rect -683 -37 -563 -21
rect -683 -71 -667 -37
rect -579 -71 -563 -37
rect -683 -118 -563 -71
rect -505 -37 -385 -21
rect -505 -71 -489 -37
rect -401 -71 -385 -37
rect -505 -118 -385 -71
rect -327 -37 -207 -21
rect -327 -71 -311 -37
rect -223 -71 -207 -37
rect -327 -118 -207 -71
rect -149 -37 -29 -21
rect -149 -71 -133 -37
rect -45 -71 -29 -37
rect -149 -118 -29 -71
rect 29 -37 149 -21
rect 29 -71 45 -37
rect 133 -71 149 -37
rect 29 -118 149 -71
rect 207 -37 327 -21
rect 207 -71 223 -37
rect 311 -71 327 -37
rect 207 -118 327 -71
rect 385 -37 505 -21
rect 385 -71 401 -37
rect 489 -71 505 -37
rect 385 -118 505 -71
rect 563 -37 683 -21
rect 563 -71 579 -37
rect 667 -71 683 -37
rect 563 -118 683 -71
rect 741 -37 861 -21
rect 741 -71 757 -37
rect 845 -71 861 -37
rect 741 -118 861 -71
rect 919 -37 1039 -21
rect 919 -71 935 -37
rect 1023 -71 1039 -37
rect 919 -118 1039 -71
rect 1097 -37 1217 -21
rect 1097 -71 1113 -37
rect 1201 -71 1217 -37
rect 1097 -118 1217 -71
rect 1275 -37 1395 -21
rect 1275 -71 1291 -37
rect 1379 -71 1395 -37
rect 1275 -118 1395 -71
rect 1453 -37 1573 -21
rect 1453 -71 1469 -37
rect 1557 -71 1573 -37
rect 1453 -118 1573 -71
rect 1631 -37 1751 -21
rect 1631 -71 1647 -37
rect 1735 -71 1751 -37
rect 1631 -118 1751 -71
rect 1809 -37 1929 -21
rect 1809 -71 1825 -37
rect 1913 -71 1929 -37
rect 1809 -118 1929 -71
rect 1987 -37 2107 -21
rect 1987 -71 2003 -37
rect 2091 -71 2107 -37
rect 1987 -118 2107 -71
rect 2165 -37 2285 -21
rect 2165 -71 2181 -37
rect 2269 -71 2285 -37
rect 2165 -118 2285 -71
rect 2343 -37 2463 -21
rect 2343 -71 2359 -37
rect 2447 -71 2463 -37
rect 2343 -118 2463 -71
rect 2521 -37 2641 -21
rect 2521 -71 2537 -37
rect 2625 -71 2641 -37
rect 2521 -118 2641 -71
rect 2699 -37 2819 -21
rect 2699 -71 2715 -37
rect 2803 -71 2819 -37
rect 2699 -118 2819 -71
rect 2877 -37 2997 -21
rect 2877 -71 2893 -37
rect 2981 -71 2997 -37
rect 2877 -118 2997 -71
rect 3055 -37 3175 -21
rect 3055 -71 3071 -37
rect 3159 -71 3175 -37
rect 3055 -118 3175 -71
rect 3233 -37 3353 -21
rect 3233 -71 3249 -37
rect 3337 -71 3353 -37
rect 3233 -118 3353 -71
rect 3411 -37 3531 -21
rect 3411 -71 3427 -37
rect 3515 -71 3531 -37
rect 3411 -118 3531 -71
rect 3589 -37 3709 -21
rect 3589 -71 3605 -37
rect 3693 -71 3709 -37
rect 3589 -118 3709 -71
rect 3767 -37 3887 -21
rect 3767 -71 3783 -37
rect 3871 -71 3887 -37
rect 3767 -118 3887 -71
rect 3945 -37 4065 -21
rect 3945 -71 3961 -37
rect 4049 -71 4065 -37
rect 3945 -118 4065 -71
rect 4123 -37 4243 -21
rect 4123 -71 4139 -37
rect 4227 -71 4243 -37
rect 4123 -118 4243 -71
rect 4301 -37 4421 -21
rect 4301 -71 4317 -37
rect 4405 -71 4421 -37
rect 4301 -118 4421 -71
rect 4479 -37 4599 -21
rect 4479 -71 4495 -37
rect 4583 -71 4599 -37
rect 4479 -118 4599 -71
rect 4657 -37 4777 -21
rect 4657 -71 4673 -37
rect 4761 -71 4777 -37
rect 4657 -118 4777 -71
rect 4835 -37 4955 -21
rect 4835 -71 4851 -37
rect 4939 -71 4955 -37
rect 4835 -118 4955 -71
rect 5013 -37 5133 -21
rect 5013 -71 5029 -37
rect 5117 -71 5133 -37
rect 5013 -118 5133 -71
rect 5191 -37 5311 -21
rect 5191 -71 5207 -37
rect 5295 -71 5311 -37
rect 5191 -118 5311 -71
rect 5369 -37 5489 -21
rect 5369 -71 5385 -37
rect 5473 -71 5489 -37
rect 5369 -118 5489 -71
rect 5547 -37 5667 -21
rect 5547 -71 5563 -37
rect 5651 -71 5667 -37
rect 5547 -118 5667 -71
rect 5725 -37 5845 -21
rect 5725 -71 5741 -37
rect 5829 -71 5845 -37
rect 5725 -118 5845 -71
rect 5903 -37 6023 -21
rect 5903 -71 5919 -37
rect 6007 -71 6023 -37
rect 5903 -118 6023 -71
rect 6081 -37 6201 -21
rect 6081 -71 6097 -37
rect 6185 -71 6201 -37
rect 6081 -118 6201 -71
rect 6259 -37 6379 -21
rect 6259 -71 6275 -37
rect 6363 -71 6379 -37
rect 6259 -118 6379 -71
rect 6437 -37 6557 -21
rect 6437 -71 6453 -37
rect 6541 -71 6557 -37
rect 6437 -118 6557 -71
rect 6615 -37 6735 -21
rect 6615 -71 6631 -37
rect 6719 -71 6735 -37
rect 6615 -118 6735 -71
rect 6793 -37 6913 -21
rect 6793 -71 6809 -37
rect 6897 -71 6913 -37
rect 6793 -118 6913 -71
rect 6971 -37 7091 -21
rect 6971 -71 6987 -37
rect 7075 -71 7091 -37
rect 6971 -118 7091 -71
rect 7149 -37 7269 -21
rect 7149 -71 7165 -37
rect 7253 -71 7269 -37
rect 7149 -118 7269 -71
rect 7327 -37 7447 -21
rect 7327 -71 7343 -37
rect 7431 -71 7447 -37
rect 7327 -118 7447 -71
rect 7505 -37 7625 -21
rect 7505 -71 7521 -37
rect 7609 -71 7625 -37
rect 7505 -118 7625 -71
rect 7683 -37 7803 -21
rect 7683 -71 7699 -37
rect 7787 -71 7803 -37
rect 7683 -118 7803 -71
rect 7861 -37 7981 -21
rect 7861 -71 7877 -37
rect 7965 -71 7981 -37
rect 7861 -118 7981 -71
rect -7981 -1365 -7861 -1318
rect -7981 -1399 -7965 -1365
rect -7877 -1399 -7861 -1365
rect -7981 -1415 -7861 -1399
rect -7803 -1365 -7683 -1318
rect -7803 -1399 -7787 -1365
rect -7699 -1399 -7683 -1365
rect -7803 -1415 -7683 -1399
rect -7625 -1365 -7505 -1318
rect -7625 -1399 -7609 -1365
rect -7521 -1399 -7505 -1365
rect -7625 -1415 -7505 -1399
rect -7447 -1365 -7327 -1318
rect -7447 -1399 -7431 -1365
rect -7343 -1399 -7327 -1365
rect -7447 -1415 -7327 -1399
rect -7269 -1365 -7149 -1318
rect -7269 -1399 -7253 -1365
rect -7165 -1399 -7149 -1365
rect -7269 -1415 -7149 -1399
rect -7091 -1365 -6971 -1318
rect -7091 -1399 -7075 -1365
rect -6987 -1399 -6971 -1365
rect -7091 -1415 -6971 -1399
rect -6913 -1365 -6793 -1318
rect -6913 -1399 -6897 -1365
rect -6809 -1399 -6793 -1365
rect -6913 -1415 -6793 -1399
rect -6735 -1365 -6615 -1318
rect -6735 -1399 -6719 -1365
rect -6631 -1399 -6615 -1365
rect -6735 -1415 -6615 -1399
rect -6557 -1365 -6437 -1318
rect -6557 -1399 -6541 -1365
rect -6453 -1399 -6437 -1365
rect -6557 -1415 -6437 -1399
rect -6379 -1365 -6259 -1318
rect -6379 -1399 -6363 -1365
rect -6275 -1399 -6259 -1365
rect -6379 -1415 -6259 -1399
rect -6201 -1365 -6081 -1318
rect -6201 -1399 -6185 -1365
rect -6097 -1399 -6081 -1365
rect -6201 -1415 -6081 -1399
rect -6023 -1365 -5903 -1318
rect -6023 -1399 -6007 -1365
rect -5919 -1399 -5903 -1365
rect -6023 -1415 -5903 -1399
rect -5845 -1365 -5725 -1318
rect -5845 -1399 -5829 -1365
rect -5741 -1399 -5725 -1365
rect -5845 -1415 -5725 -1399
rect -5667 -1365 -5547 -1318
rect -5667 -1399 -5651 -1365
rect -5563 -1399 -5547 -1365
rect -5667 -1415 -5547 -1399
rect -5489 -1365 -5369 -1318
rect -5489 -1399 -5473 -1365
rect -5385 -1399 -5369 -1365
rect -5489 -1415 -5369 -1399
rect -5311 -1365 -5191 -1318
rect -5311 -1399 -5295 -1365
rect -5207 -1399 -5191 -1365
rect -5311 -1415 -5191 -1399
rect -5133 -1365 -5013 -1318
rect -5133 -1399 -5117 -1365
rect -5029 -1399 -5013 -1365
rect -5133 -1415 -5013 -1399
rect -4955 -1365 -4835 -1318
rect -4955 -1399 -4939 -1365
rect -4851 -1399 -4835 -1365
rect -4955 -1415 -4835 -1399
rect -4777 -1365 -4657 -1318
rect -4777 -1399 -4761 -1365
rect -4673 -1399 -4657 -1365
rect -4777 -1415 -4657 -1399
rect -4599 -1365 -4479 -1318
rect -4599 -1399 -4583 -1365
rect -4495 -1399 -4479 -1365
rect -4599 -1415 -4479 -1399
rect -4421 -1365 -4301 -1318
rect -4421 -1399 -4405 -1365
rect -4317 -1399 -4301 -1365
rect -4421 -1415 -4301 -1399
rect -4243 -1365 -4123 -1318
rect -4243 -1399 -4227 -1365
rect -4139 -1399 -4123 -1365
rect -4243 -1415 -4123 -1399
rect -4065 -1365 -3945 -1318
rect -4065 -1399 -4049 -1365
rect -3961 -1399 -3945 -1365
rect -4065 -1415 -3945 -1399
rect -3887 -1365 -3767 -1318
rect -3887 -1399 -3871 -1365
rect -3783 -1399 -3767 -1365
rect -3887 -1415 -3767 -1399
rect -3709 -1365 -3589 -1318
rect -3709 -1399 -3693 -1365
rect -3605 -1399 -3589 -1365
rect -3709 -1415 -3589 -1399
rect -3531 -1365 -3411 -1318
rect -3531 -1399 -3515 -1365
rect -3427 -1399 -3411 -1365
rect -3531 -1415 -3411 -1399
rect -3353 -1365 -3233 -1318
rect -3353 -1399 -3337 -1365
rect -3249 -1399 -3233 -1365
rect -3353 -1415 -3233 -1399
rect -3175 -1365 -3055 -1318
rect -3175 -1399 -3159 -1365
rect -3071 -1399 -3055 -1365
rect -3175 -1415 -3055 -1399
rect -2997 -1365 -2877 -1318
rect -2997 -1399 -2981 -1365
rect -2893 -1399 -2877 -1365
rect -2997 -1415 -2877 -1399
rect -2819 -1365 -2699 -1318
rect -2819 -1399 -2803 -1365
rect -2715 -1399 -2699 -1365
rect -2819 -1415 -2699 -1399
rect -2641 -1365 -2521 -1318
rect -2641 -1399 -2625 -1365
rect -2537 -1399 -2521 -1365
rect -2641 -1415 -2521 -1399
rect -2463 -1365 -2343 -1318
rect -2463 -1399 -2447 -1365
rect -2359 -1399 -2343 -1365
rect -2463 -1415 -2343 -1399
rect -2285 -1365 -2165 -1318
rect -2285 -1399 -2269 -1365
rect -2181 -1399 -2165 -1365
rect -2285 -1415 -2165 -1399
rect -2107 -1365 -1987 -1318
rect -2107 -1399 -2091 -1365
rect -2003 -1399 -1987 -1365
rect -2107 -1415 -1987 -1399
rect -1929 -1365 -1809 -1318
rect -1929 -1399 -1913 -1365
rect -1825 -1399 -1809 -1365
rect -1929 -1415 -1809 -1399
rect -1751 -1365 -1631 -1318
rect -1751 -1399 -1735 -1365
rect -1647 -1399 -1631 -1365
rect -1751 -1415 -1631 -1399
rect -1573 -1365 -1453 -1318
rect -1573 -1399 -1557 -1365
rect -1469 -1399 -1453 -1365
rect -1573 -1415 -1453 -1399
rect -1395 -1365 -1275 -1318
rect -1395 -1399 -1379 -1365
rect -1291 -1399 -1275 -1365
rect -1395 -1415 -1275 -1399
rect -1217 -1365 -1097 -1318
rect -1217 -1399 -1201 -1365
rect -1113 -1399 -1097 -1365
rect -1217 -1415 -1097 -1399
rect -1039 -1365 -919 -1318
rect -1039 -1399 -1023 -1365
rect -935 -1399 -919 -1365
rect -1039 -1415 -919 -1399
rect -861 -1365 -741 -1318
rect -861 -1399 -845 -1365
rect -757 -1399 -741 -1365
rect -861 -1415 -741 -1399
rect -683 -1365 -563 -1318
rect -683 -1399 -667 -1365
rect -579 -1399 -563 -1365
rect -683 -1415 -563 -1399
rect -505 -1365 -385 -1318
rect -505 -1399 -489 -1365
rect -401 -1399 -385 -1365
rect -505 -1415 -385 -1399
rect -327 -1365 -207 -1318
rect -327 -1399 -311 -1365
rect -223 -1399 -207 -1365
rect -327 -1415 -207 -1399
rect -149 -1365 -29 -1318
rect -149 -1399 -133 -1365
rect -45 -1399 -29 -1365
rect -149 -1415 -29 -1399
rect 29 -1365 149 -1318
rect 29 -1399 45 -1365
rect 133 -1399 149 -1365
rect 29 -1415 149 -1399
rect 207 -1365 327 -1318
rect 207 -1399 223 -1365
rect 311 -1399 327 -1365
rect 207 -1415 327 -1399
rect 385 -1365 505 -1318
rect 385 -1399 401 -1365
rect 489 -1399 505 -1365
rect 385 -1415 505 -1399
rect 563 -1365 683 -1318
rect 563 -1399 579 -1365
rect 667 -1399 683 -1365
rect 563 -1415 683 -1399
rect 741 -1365 861 -1318
rect 741 -1399 757 -1365
rect 845 -1399 861 -1365
rect 741 -1415 861 -1399
rect 919 -1365 1039 -1318
rect 919 -1399 935 -1365
rect 1023 -1399 1039 -1365
rect 919 -1415 1039 -1399
rect 1097 -1365 1217 -1318
rect 1097 -1399 1113 -1365
rect 1201 -1399 1217 -1365
rect 1097 -1415 1217 -1399
rect 1275 -1365 1395 -1318
rect 1275 -1399 1291 -1365
rect 1379 -1399 1395 -1365
rect 1275 -1415 1395 -1399
rect 1453 -1365 1573 -1318
rect 1453 -1399 1469 -1365
rect 1557 -1399 1573 -1365
rect 1453 -1415 1573 -1399
rect 1631 -1365 1751 -1318
rect 1631 -1399 1647 -1365
rect 1735 -1399 1751 -1365
rect 1631 -1415 1751 -1399
rect 1809 -1365 1929 -1318
rect 1809 -1399 1825 -1365
rect 1913 -1399 1929 -1365
rect 1809 -1415 1929 -1399
rect 1987 -1365 2107 -1318
rect 1987 -1399 2003 -1365
rect 2091 -1399 2107 -1365
rect 1987 -1415 2107 -1399
rect 2165 -1365 2285 -1318
rect 2165 -1399 2181 -1365
rect 2269 -1399 2285 -1365
rect 2165 -1415 2285 -1399
rect 2343 -1365 2463 -1318
rect 2343 -1399 2359 -1365
rect 2447 -1399 2463 -1365
rect 2343 -1415 2463 -1399
rect 2521 -1365 2641 -1318
rect 2521 -1399 2537 -1365
rect 2625 -1399 2641 -1365
rect 2521 -1415 2641 -1399
rect 2699 -1365 2819 -1318
rect 2699 -1399 2715 -1365
rect 2803 -1399 2819 -1365
rect 2699 -1415 2819 -1399
rect 2877 -1365 2997 -1318
rect 2877 -1399 2893 -1365
rect 2981 -1399 2997 -1365
rect 2877 -1415 2997 -1399
rect 3055 -1365 3175 -1318
rect 3055 -1399 3071 -1365
rect 3159 -1399 3175 -1365
rect 3055 -1415 3175 -1399
rect 3233 -1365 3353 -1318
rect 3233 -1399 3249 -1365
rect 3337 -1399 3353 -1365
rect 3233 -1415 3353 -1399
rect 3411 -1365 3531 -1318
rect 3411 -1399 3427 -1365
rect 3515 -1399 3531 -1365
rect 3411 -1415 3531 -1399
rect 3589 -1365 3709 -1318
rect 3589 -1399 3605 -1365
rect 3693 -1399 3709 -1365
rect 3589 -1415 3709 -1399
rect 3767 -1365 3887 -1318
rect 3767 -1399 3783 -1365
rect 3871 -1399 3887 -1365
rect 3767 -1415 3887 -1399
rect 3945 -1365 4065 -1318
rect 3945 -1399 3961 -1365
rect 4049 -1399 4065 -1365
rect 3945 -1415 4065 -1399
rect 4123 -1365 4243 -1318
rect 4123 -1399 4139 -1365
rect 4227 -1399 4243 -1365
rect 4123 -1415 4243 -1399
rect 4301 -1365 4421 -1318
rect 4301 -1399 4317 -1365
rect 4405 -1399 4421 -1365
rect 4301 -1415 4421 -1399
rect 4479 -1365 4599 -1318
rect 4479 -1399 4495 -1365
rect 4583 -1399 4599 -1365
rect 4479 -1415 4599 -1399
rect 4657 -1365 4777 -1318
rect 4657 -1399 4673 -1365
rect 4761 -1399 4777 -1365
rect 4657 -1415 4777 -1399
rect 4835 -1365 4955 -1318
rect 4835 -1399 4851 -1365
rect 4939 -1399 4955 -1365
rect 4835 -1415 4955 -1399
rect 5013 -1365 5133 -1318
rect 5013 -1399 5029 -1365
rect 5117 -1399 5133 -1365
rect 5013 -1415 5133 -1399
rect 5191 -1365 5311 -1318
rect 5191 -1399 5207 -1365
rect 5295 -1399 5311 -1365
rect 5191 -1415 5311 -1399
rect 5369 -1365 5489 -1318
rect 5369 -1399 5385 -1365
rect 5473 -1399 5489 -1365
rect 5369 -1415 5489 -1399
rect 5547 -1365 5667 -1318
rect 5547 -1399 5563 -1365
rect 5651 -1399 5667 -1365
rect 5547 -1415 5667 -1399
rect 5725 -1365 5845 -1318
rect 5725 -1399 5741 -1365
rect 5829 -1399 5845 -1365
rect 5725 -1415 5845 -1399
rect 5903 -1365 6023 -1318
rect 5903 -1399 5919 -1365
rect 6007 -1399 6023 -1365
rect 5903 -1415 6023 -1399
rect 6081 -1365 6201 -1318
rect 6081 -1399 6097 -1365
rect 6185 -1399 6201 -1365
rect 6081 -1415 6201 -1399
rect 6259 -1365 6379 -1318
rect 6259 -1399 6275 -1365
rect 6363 -1399 6379 -1365
rect 6259 -1415 6379 -1399
rect 6437 -1365 6557 -1318
rect 6437 -1399 6453 -1365
rect 6541 -1399 6557 -1365
rect 6437 -1415 6557 -1399
rect 6615 -1365 6735 -1318
rect 6615 -1399 6631 -1365
rect 6719 -1399 6735 -1365
rect 6615 -1415 6735 -1399
rect 6793 -1365 6913 -1318
rect 6793 -1399 6809 -1365
rect 6897 -1399 6913 -1365
rect 6793 -1415 6913 -1399
rect 6971 -1365 7091 -1318
rect 6971 -1399 6987 -1365
rect 7075 -1399 7091 -1365
rect 6971 -1415 7091 -1399
rect 7149 -1365 7269 -1318
rect 7149 -1399 7165 -1365
rect 7253 -1399 7269 -1365
rect 7149 -1415 7269 -1399
rect 7327 -1365 7447 -1318
rect 7327 -1399 7343 -1365
rect 7431 -1399 7447 -1365
rect 7327 -1415 7447 -1399
rect 7505 -1365 7625 -1318
rect 7505 -1399 7521 -1365
rect 7609 -1399 7625 -1365
rect 7505 -1415 7625 -1399
rect 7683 -1365 7803 -1318
rect 7683 -1399 7699 -1365
rect 7787 -1399 7803 -1365
rect 7683 -1415 7803 -1399
rect 7861 -1365 7981 -1318
rect 7861 -1399 7877 -1365
rect 7965 -1399 7981 -1365
rect 7861 -1415 7981 -1399
<< polycont >>
rect -7965 1365 -7877 1399
rect -7787 1365 -7699 1399
rect -7609 1365 -7521 1399
rect -7431 1365 -7343 1399
rect -7253 1365 -7165 1399
rect -7075 1365 -6987 1399
rect -6897 1365 -6809 1399
rect -6719 1365 -6631 1399
rect -6541 1365 -6453 1399
rect -6363 1365 -6275 1399
rect -6185 1365 -6097 1399
rect -6007 1365 -5919 1399
rect -5829 1365 -5741 1399
rect -5651 1365 -5563 1399
rect -5473 1365 -5385 1399
rect -5295 1365 -5207 1399
rect -5117 1365 -5029 1399
rect -4939 1365 -4851 1399
rect -4761 1365 -4673 1399
rect -4583 1365 -4495 1399
rect -4405 1365 -4317 1399
rect -4227 1365 -4139 1399
rect -4049 1365 -3961 1399
rect -3871 1365 -3783 1399
rect -3693 1365 -3605 1399
rect -3515 1365 -3427 1399
rect -3337 1365 -3249 1399
rect -3159 1365 -3071 1399
rect -2981 1365 -2893 1399
rect -2803 1365 -2715 1399
rect -2625 1365 -2537 1399
rect -2447 1365 -2359 1399
rect -2269 1365 -2181 1399
rect -2091 1365 -2003 1399
rect -1913 1365 -1825 1399
rect -1735 1365 -1647 1399
rect -1557 1365 -1469 1399
rect -1379 1365 -1291 1399
rect -1201 1365 -1113 1399
rect -1023 1365 -935 1399
rect -845 1365 -757 1399
rect -667 1365 -579 1399
rect -489 1365 -401 1399
rect -311 1365 -223 1399
rect -133 1365 -45 1399
rect 45 1365 133 1399
rect 223 1365 311 1399
rect 401 1365 489 1399
rect 579 1365 667 1399
rect 757 1365 845 1399
rect 935 1365 1023 1399
rect 1113 1365 1201 1399
rect 1291 1365 1379 1399
rect 1469 1365 1557 1399
rect 1647 1365 1735 1399
rect 1825 1365 1913 1399
rect 2003 1365 2091 1399
rect 2181 1365 2269 1399
rect 2359 1365 2447 1399
rect 2537 1365 2625 1399
rect 2715 1365 2803 1399
rect 2893 1365 2981 1399
rect 3071 1365 3159 1399
rect 3249 1365 3337 1399
rect 3427 1365 3515 1399
rect 3605 1365 3693 1399
rect 3783 1365 3871 1399
rect 3961 1365 4049 1399
rect 4139 1365 4227 1399
rect 4317 1365 4405 1399
rect 4495 1365 4583 1399
rect 4673 1365 4761 1399
rect 4851 1365 4939 1399
rect 5029 1365 5117 1399
rect 5207 1365 5295 1399
rect 5385 1365 5473 1399
rect 5563 1365 5651 1399
rect 5741 1365 5829 1399
rect 5919 1365 6007 1399
rect 6097 1365 6185 1399
rect 6275 1365 6363 1399
rect 6453 1365 6541 1399
rect 6631 1365 6719 1399
rect 6809 1365 6897 1399
rect 6987 1365 7075 1399
rect 7165 1365 7253 1399
rect 7343 1365 7431 1399
rect 7521 1365 7609 1399
rect 7699 1365 7787 1399
rect 7877 1365 7965 1399
rect -7965 37 -7877 71
rect -7787 37 -7699 71
rect -7609 37 -7521 71
rect -7431 37 -7343 71
rect -7253 37 -7165 71
rect -7075 37 -6987 71
rect -6897 37 -6809 71
rect -6719 37 -6631 71
rect -6541 37 -6453 71
rect -6363 37 -6275 71
rect -6185 37 -6097 71
rect -6007 37 -5919 71
rect -5829 37 -5741 71
rect -5651 37 -5563 71
rect -5473 37 -5385 71
rect -5295 37 -5207 71
rect -5117 37 -5029 71
rect -4939 37 -4851 71
rect -4761 37 -4673 71
rect -4583 37 -4495 71
rect -4405 37 -4317 71
rect -4227 37 -4139 71
rect -4049 37 -3961 71
rect -3871 37 -3783 71
rect -3693 37 -3605 71
rect -3515 37 -3427 71
rect -3337 37 -3249 71
rect -3159 37 -3071 71
rect -2981 37 -2893 71
rect -2803 37 -2715 71
rect -2625 37 -2537 71
rect -2447 37 -2359 71
rect -2269 37 -2181 71
rect -2091 37 -2003 71
rect -1913 37 -1825 71
rect -1735 37 -1647 71
rect -1557 37 -1469 71
rect -1379 37 -1291 71
rect -1201 37 -1113 71
rect -1023 37 -935 71
rect -845 37 -757 71
rect -667 37 -579 71
rect -489 37 -401 71
rect -311 37 -223 71
rect -133 37 -45 71
rect 45 37 133 71
rect 223 37 311 71
rect 401 37 489 71
rect 579 37 667 71
rect 757 37 845 71
rect 935 37 1023 71
rect 1113 37 1201 71
rect 1291 37 1379 71
rect 1469 37 1557 71
rect 1647 37 1735 71
rect 1825 37 1913 71
rect 2003 37 2091 71
rect 2181 37 2269 71
rect 2359 37 2447 71
rect 2537 37 2625 71
rect 2715 37 2803 71
rect 2893 37 2981 71
rect 3071 37 3159 71
rect 3249 37 3337 71
rect 3427 37 3515 71
rect 3605 37 3693 71
rect 3783 37 3871 71
rect 3961 37 4049 71
rect 4139 37 4227 71
rect 4317 37 4405 71
rect 4495 37 4583 71
rect 4673 37 4761 71
rect 4851 37 4939 71
rect 5029 37 5117 71
rect 5207 37 5295 71
rect 5385 37 5473 71
rect 5563 37 5651 71
rect 5741 37 5829 71
rect 5919 37 6007 71
rect 6097 37 6185 71
rect 6275 37 6363 71
rect 6453 37 6541 71
rect 6631 37 6719 71
rect 6809 37 6897 71
rect 6987 37 7075 71
rect 7165 37 7253 71
rect 7343 37 7431 71
rect 7521 37 7609 71
rect 7699 37 7787 71
rect 7877 37 7965 71
rect -7965 -71 -7877 -37
rect -7787 -71 -7699 -37
rect -7609 -71 -7521 -37
rect -7431 -71 -7343 -37
rect -7253 -71 -7165 -37
rect -7075 -71 -6987 -37
rect -6897 -71 -6809 -37
rect -6719 -71 -6631 -37
rect -6541 -71 -6453 -37
rect -6363 -71 -6275 -37
rect -6185 -71 -6097 -37
rect -6007 -71 -5919 -37
rect -5829 -71 -5741 -37
rect -5651 -71 -5563 -37
rect -5473 -71 -5385 -37
rect -5295 -71 -5207 -37
rect -5117 -71 -5029 -37
rect -4939 -71 -4851 -37
rect -4761 -71 -4673 -37
rect -4583 -71 -4495 -37
rect -4405 -71 -4317 -37
rect -4227 -71 -4139 -37
rect -4049 -71 -3961 -37
rect -3871 -71 -3783 -37
rect -3693 -71 -3605 -37
rect -3515 -71 -3427 -37
rect -3337 -71 -3249 -37
rect -3159 -71 -3071 -37
rect -2981 -71 -2893 -37
rect -2803 -71 -2715 -37
rect -2625 -71 -2537 -37
rect -2447 -71 -2359 -37
rect -2269 -71 -2181 -37
rect -2091 -71 -2003 -37
rect -1913 -71 -1825 -37
rect -1735 -71 -1647 -37
rect -1557 -71 -1469 -37
rect -1379 -71 -1291 -37
rect -1201 -71 -1113 -37
rect -1023 -71 -935 -37
rect -845 -71 -757 -37
rect -667 -71 -579 -37
rect -489 -71 -401 -37
rect -311 -71 -223 -37
rect -133 -71 -45 -37
rect 45 -71 133 -37
rect 223 -71 311 -37
rect 401 -71 489 -37
rect 579 -71 667 -37
rect 757 -71 845 -37
rect 935 -71 1023 -37
rect 1113 -71 1201 -37
rect 1291 -71 1379 -37
rect 1469 -71 1557 -37
rect 1647 -71 1735 -37
rect 1825 -71 1913 -37
rect 2003 -71 2091 -37
rect 2181 -71 2269 -37
rect 2359 -71 2447 -37
rect 2537 -71 2625 -37
rect 2715 -71 2803 -37
rect 2893 -71 2981 -37
rect 3071 -71 3159 -37
rect 3249 -71 3337 -37
rect 3427 -71 3515 -37
rect 3605 -71 3693 -37
rect 3783 -71 3871 -37
rect 3961 -71 4049 -37
rect 4139 -71 4227 -37
rect 4317 -71 4405 -37
rect 4495 -71 4583 -37
rect 4673 -71 4761 -37
rect 4851 -71 4939 -37
rect 5029 -71 5117 -37
rect 5207 -71 5295 -37
rect 5385 -71 5473 -37
rect 5563 -71 5651 -37
rect 5741 -71 5829 -37
rect 5919 -71 6007 -37
rect 6097 -71 6185 -37
rect 6275 -71 6363 -37
rect 6453 -71 6541 -37
rect 6631 -71 6719 -37
rect 6809 -71 6897 -37
rect 6987 -71 7075 -37
rect 7165 -71 7253 -37
rect 7343 -71 7431 -37
rect 7521 -71 7609 -37
rect 7699 -71 7787 -37
rect 7877 -71 7965 -37
rect -7965 -1399 -7877 -1365
rect -7787 -1399 -7699 -1365
rect -7609 -1399 -7521 -1365
rect -7431 -1399 -7343 -1365
rect -7253 -1399 -7165 -1365
rect -7075 -1399 -6987 -1365
rect -6897 -1399 -6809 -1365
rect -6719 -1399 -6631 -1365
rect -6541 -1399 -6453 -1365
rect -6363 -1399 -6275 -1365
rect -6185 -1399 -6097 -1365
rect -6007 -1399 -5919 -1365
rect -5829 -1399 -5741 -1365
rect -5651 -1399 -5563 -1365
rect -5473 -1399 -5385 -1365
rect -5295 -1399 -5207 -1365
rect -5117 -1399 -5029 -1365
rect -4939 -1399 -4851 -1365
rect -4761 -1399 -4673 -1365
rect -4583 -1399 -4495 -1365
rect -4405 -1399 -4317 -1365
rect -4227 -1399 -4139 -1365
rect -4049 -1399 -3961 -1365
rect -3871 -1399 -3783 -1365
rect -3693 -1399 -3605 -1365
rect -3515 -1399 -3427 -1365
rect -3337 -1399 -3249 -1365
rect -3159 -1399 -3071 -1365
rect -2981 -1399 -2893 -1365
rect -2803 -1399 -2715 -1365
rect -2625 -1399 -2537 -1365
rect -2447 -1399 -2359 -1365
rect -2269 -1399 -2181 -1365
rect -2091 -1399 -2003 -1365
rect -1913 -1399 -1825 -1365
rect -1735 -1399 -1647 -1365
rect -1557 -1399 -1469 -1365
rect -1379 -1399 -1291 -1365
rect -1201 -1399 -1113 -1365
rect -1023 -1399 -935 -1365
rect -845 -1399 -757 -1365
rect -667 -1399 -579 -1365
rect -489 -1399 -401 -1365
rect -311 -1399 -223 -1365
rect -133 -1399 -45 -1365
rect 45 -1399 133 -1365
rect 223 -1399 311 -1365
rect 401 -1399 489 -1365
rect 579 -1399 667 -1365
rect 757 -1399 845 -1365
rect 935 -1399 1023 -1365
rect 1113 -1399 1201 -1365
rect 1291 -1399 1379 -1365
rect 1469 -1399 1557 -1365
rect 1647 -1399 1735 -1365
rect 1825 -1399 1913 -1365
rect 2003 -1399 2091 -1365
rect 2181 -1399 2269 -1365
rect 2359 -1399 2447 -1365
rect 2537 -1399 2625 -1365
rect 2715 -1399 2803 -1365
rect 2893 -1399 2981 -1365
rect 3071 -1399 3159 -1365
rect 3249 -1399 3337 -1365
rect 3427 -1399 3515 -1365
rect 3605 -1399 3693 -1365
rect 3783 -1399 3871 -1365
rect 3961 -1399 4049 -1365
rect 4139 -1399 4227 -1365
rect 4317 -1399 4405 -1365
rect 4495 -1399 4583 -1365
rect 4673 -1399 4761 -1365
rect 4851 -1399 4939 -1365
rect 5029 -1399 5117 -1365
rect 5207 -1399 5295 -1365
rect 5385 -1399 5473 -1365
rect 5563 -1399 5651 -1365
rect 5741 -1399 5829 -1365
rect 5919 -1399 6007 -1365
rect 6097 -1399 6185 -1365
rect 6275 -1399 6363 -1365
rect 6453 -1399 6541 -1365
rect 6631 -1399 6719 -1365
rect 6809 -1399 6897 -1365
rect 6987 -1399 7075 -1365
rect 7165 -1399 7253 -1365
rect 7343 -1399 7431 -1365
rect 7521 -1399 7609 -1365
rect 7699 -1399 7787 -1365
rect 7877 -1399 7965 -1365
<< locali >>
rect -8141 1467 -8045 1501
rect 8045 1467 8141 1501
rect -8141 1405 -8107 1467
rect 8107 1405 8141 1467
rect -7981 1365 -7965 1399
rect -7877 1365 -7861 1399
rect -7803 1365 -7787 1399
rect -7699 1365 -7683 1399
rect -7625 1365 -7609 1399
rect -7521 1365 -7505 1399
rect -7447 1365 -7431 1399
rect -7343 1365 -7327 1399
rect -7269 1365 -7253 1399
rect -7165 1365 -7149 1399
rect -7091 1365 -7075 1399
rect -6987 1365 -6971 1399
rect -6913 1365 -6897 1399
rect -6809 1365 -6793 1399
rect -6735 1365 -6719 1399
rect -6631 1365 -6615 1399
rect -6557 1365 -6541 1399
rect -6453 1365 -6437 1399
rect -6379 1365 -6363 1399
rect -6275 1365 -6259 1399
rect -6201 1365 -6185 1399
rect -6097 1365 -6081 1399
rect -6023 1365 -6007 1399
rect -5919 1365 -5903 1399
rect -5845 1365 -5829 1399
rect -5741 1365 -5725 1399
rect -5667 1365 -5651 1399
rect -5563 1365 -5547 1399
rect -5489 1365 -5473 1399
rect -5385 1365 -5369 1399
rect -5311 1365 -5295 1399
rect -5207 1365 -5191 1399
rect -5133 1365 -5117 1399
rect -5029 1365 -5013 1399
rect -4955 1365 -4939 1399
rect -4851 1365 -4835 1399
rect -4777 1365 -4761 1399
rect -4673 1365 -4657 1399
rect -4599 1365 -4583 1399
rect -4495 1365 -4479 1399
rect -4421 1365 -4405 1399
rect -4317 1365 -4301 1399
rect -4243 1365 -4227 1399
rect -4139 1365 -4123 1399
rect -4065 1365 -4049 1399
rect -3961 1365 -3945 1399
rect -3887 1365 -3871 1399
rect -3783 1365 -3767 1399
rect -3709 1365 -3693 1399
rect -3605 1365 -3589 1399
rect -3531 1365 -3515 1399
rect -3427 1365 -3411 1399
rect -3353 1365 -3337 1399
rect -3249 1365 -3233 1399
rect -3175 1365 -3159 1399
rect -3071 1365 -3055 1399
rect -2997 1365 -2981 1399
rect -2893 1365 -2877 1399
rect -2819 1365 -2803 1399
rect -2715 1365 -2699 1399
rect -2641 1365 -2625 1399
rect -2537 1365 -2521 1399
rect -2463 1365 -2447 1399
rect -2359 1365 -2343 1399
rect -2285 1365 -2269 1399
rect -2181 1365 -2165 1399
rect -2107 1365 -2091 1399
rect -2003 1365 -1987 1399
rect -1929 1365 -1913 1399
rect -1825 1365 -1809 1399
rect -1751 1365 -1735 1399
rect -1647 1365 -1631 1399
rect -1573 1365 -1557 1399
rect -1469 1365 -1453 1399
rect -1395 1365 -1379 1399
rect -1291 1365 -1275 1399
rect -1217 1365 -1201 1399
rect -1113 1365 -1097 1399
rect -1039 1365 -1023 1399
rect -935 1365 -919 1399
rect -861 1365 -845 1399
rect -757 1365 -741 1399
rect -683 1365 -667 1399
rect -579 1365 -563 1399
rect -505 1365 -489 1399
rect -401 1365 -385 1399
rect -327 1365 -311 1399
rect -223 1365 -207 1399
rect -149 1365 -133 1399
rect -45 1365 -29 1399
rect 29 1365 45 1399
rect 133 1365 149 1399
rect 207 1365 223 1399
rect 311 1365 327 1399
rect 385 1365 401 1399
rect 489 1365 505 1399
rect 563 1365 579 1399
rect 667 1365 683 1399
rect 741 1365 757 1399
rect 845 1365 861 1399
rect 919 1365 935 1399
rect 1023 1365 1039 1399
rect 1097 1365 1113 1399
rect 1201 1365 1217 1399
rect 1275 1365 1291 1399
rect 1379 1365 1395 1399
rect 1453 1365 1469 1399
rect 1557 1365 1573 1399
rect 1631 1365 1647 1399
rect 1735 1365 1751 1399
rect 1809 1365 1825 1399
rect 1913 1365 1929 1399
rect 1987 1365 2003 1399
rect 2091 1365 2107 1399
rect 2165 1365 2181 1399
rect 2269 1365 2285 1399
rect 2343 1365 2359 1399
rect 2447 1365 2463 1399
rect 2521 1365 2537 1399
rect 2625 1365 2641 1399
rect 2699 1365 2715 1399
rect 2803 1365 2819 1399
rect 2877 1365 2893 1399
rect 2981 1365 2997 1399
rect 3055 1365 3071 1399
rect 3159 1365 3175 1399
rect 3233 1365 3249 1399
rect 3337 1365 3353 1399
rect 3411 1365 3427 1399
rect 3515 1365 3531 1399
rect 3589 1365 3605 1399
rect 3693 1365 3709 1399
rect 3767 1365 3783 1399
rect 3871 1365 3887 1399
rect 3945 1365 3961 1399
rect 4049 1365 4065 1399
rect 4123 1365 4139 1399
rect 4227 1365 4243 1399
rect 4301 1365 4317 1399
rect 4405 1365 4421 1399
rect 4479 1365 4495 1399
rect 4583 1365 4599 1399
rect 4657 1365 4673 1399
rect 4761 1365 4777 1399
rect 4835 1365 4851 1399
rect 4939 1365 4955 1399
rect 5013 1365 5029 1399
rect 5117 1365 5133 1399
rect 5191 1365 5207 1399
rect 5295 1365 5311 1399
rect 5369 1365 5385 1399
rect 5473 1365 5489 1399
rect 5547 1365 5563 1399
rect 5651 1365 5667 1399
rect 5725 1365 5741 1399
rect 5829 1365 5845 1399
rect 5903 1365 5919 1399
rect 6007 1365 6023 1399
rect 6081 1365 6097 1399
rect 6185 1365 6201 1399
rect 6259 1365 6275 1399
rect 6363 1365 6379 1399
rect 6437 1365 6453 1399
rect 6541 1365 6557 1399
rect 6615 1365 6631 1399
rect 6719 1365 6735 1399
rect 6793 1365 6809 1399
rect 6897 1365 6913 1399
rect 6971 1365 6987 1399
rect 7075 1365 7091 1399
rect 7149 1365 7165 1399
rect 7253 1365 7269 1399
rect 7327 1365 7343 1399
rect 7431 1365 7447 1399
rect 7505 1365 7521 1399
rect 7609 1365 7625 1399
rect 7683 1365 7699 1399
rect 7787 1365 7803 1399
rect 7861 1365 7877 1399
rect 7965 1365 7981 1399
rect -8027 1306 -7993 1322
rect -8027 114 -7993 130
rect -7849 1306 -7815 1322
rect -7849 114 -7815 130
rect -7671 1306 -7637 1322
rect -7671 114 -7637 130
rect -7493 1306 -7459 1322
rect -7493 114 -7459 130
rect -7315 1306 -7281 1322
rect -7315 114 -7281 130
rect -7137 1306 -7103 1322
rect -7137 114 -7103 130
rect -6959 1306 -6925 1322
rect -6959 114 -6925 130
rect -6781 1306 -6747 1322
rect -6781 114 -6747 130
rect -6603 1306 -6569 1322
rect -6603 114 -6569 130
rect -6425 1306 -6391 1322
rect -6425 114 -6391 130
rect -6247 1306 -6213 1322
rect -6247 114 -6213 130
rect -6069 1306 -6035 1322
rect -6069 114 -6035 130
rect -5891 1306 -5857 1322
rect -5891 114 -5857 130
rect -5713 1306 -5679 1322
rect -5713 114 -5679 130
rect -5535 1306 -5501 1322
rect -5535 114 -5501 130
rect -5357 1306 -5323 1322
rect -5357 114 -5323 130
rect -5179 1306 -5145 1322
rect -5179 114 -5145 130
rect -5001 1306 -4967 1322
rect -5001 114 -4967 130
rect -4823 1306 -4789 1322
rect -4823 114 -4789 130
rect -4645 1306 -4611 1322
rect -4645 114 -4611 130
rect -4467 1306 -4433 1322
rect -4467 114 -4433 130
rect -4289 1306 -4255 1322
rect -4289 114 -4255 130
rect -4111 1306 -4077 1322
rect -4111 114 -4077 130
rect -3933 1306 -3899 1322
rect -3933 114 -3899 130
rect -3755 1306 -3721 1322
rect -3755 114 -3721 130
rect -3577 1306 -3543 1322
rect -3577 114 -3543 130
rect -3399 1306 -3365 1322
rect -3399 114 -3365 130
rect -3221 1306 -3187 1322
rect -3221 114 -3187 130
rect -3043 1306 -3009 1322
rect -3043 114 -3009 130
rect -2865 1306 -2831 1322
rect -2865 114 -2831 130
rect -2687 1306 -2653 1322
rect -2687 114 -2653 130
rect -2509 1306 -2475 1322
rect -2509 114 -2475 130
rect -2331 1306 -2297 1322
rect -2331 114 -2297 130
rect -2153 1306 -2119 1322
rect -2153 114 -2119 130
rect -1975 1306 -1941 1322
rect -1975 114 -1941 130
rect -1797 1306 -1763 1322
rect -1797 114 -1763 130
rect -1619 1306 -1585 1322
rect -1619 114 -1585 130
rect -1441 1306 -1407 1322
rect -1441 114 -1407 130
rect -1263 1306 -1229 1322
rect -1263 114 -1229 130
rect -1085 1306 -1051 1322
rect -1085 114 -1051 130
rect -907 1306 -873 1322
rect -907 114 -873 130
rect -729 1306 -695 1322
rect -729 114 -695 130
rect -551 1306 -517 1322
rect -551 114 -517 130
rect -373 1306 -339 1322
rect -373 114 -339 130
rect -195 1306 -161 1322
rect -195 114 -161 130
rect -17 1306 17 1322
rect -17 114 17 130
rect 161 1306 195 1322
rect 161 114 195 130
rect 339 1306 373 1322
rect 339 114 373 130
rect 517 1306 551 1322
rect 517 114 551 130
rect 695 1306 729 1322
rect 695 114 729 130
rect 873 1306 907 1322
rect 873 114 907 130
rect 1051 1306 1085 1322
rect 1051 114 1085 130
rect 1229 1306 1263 1322
rect 1229 114 1263 130
rect 1407 1306 1441 1322
rect 1407 114 1441 130
rect 1585 1306 1619 1322
rect 1585 114 1619 130
rect 1763 1306 1797 1322
rect 1763 114 1797 130
rect 1941 1306 1975 1322
rect 1941 114 1975 130
rect 2119 1306 2153 1322
rect 2119 114 2153 130
rect 2297 1306 2331 1322
rect 2297 114 2331 130
rect 2475 1306 2509 1322
rect 2475 114 2509 130
rect 2653 1306 2687 1322
rect 2653 114 2687 130
rect 2831 1306 2865 1322
rect 2831 114 2865 130
rect 3009 1306 3043 1322
rect 3009 114 3043 130
rect 3187 1306 3221 1322
rect 3187 114 3221 130
rect 3365 1306 3399 1322
rect 3365 114 3399 130
rect 3543 1306 3577 1322
rect 3543 114 3577 130
rect 3721 1306 3755 1322
rect 3721 114 3755 130
rect 3899 1306 3933 1322
rect 3899 114 3933 130
rect 4077 1306 4111 1322
rect 4077 114 4111 130
rect 4255 1306 4289 1322
rect 4255 114 4289 130
rect 4433 1306 4467 1322
rect 4433 114 4467 130
rect 4611 1306 4645 1322
rect 4611 114 4645 130
rect 4789 1306 4823 1322
rect 4789 114 4823 130
rect 4967 1306 5001 1322
rect 4967 114 5001 130
rect 5145 1306 5179 1322
rect 5145 114 5179 130
rect 5323 1306 5357 1322
rect 5323 114 5357 130
rect 5501 1306 5535 1322
rect 5501 114 5535 130
rect 5679 1306 5713 1322
rect 5679 114 5713 130
rect 5857 1306 5891 1322
rect 5857 114 5891 130
rect 6035 1306 6069 1322
rect 6035 114 6069 130
rect 6213 1306 6247 1322
rect 6213 114 6247 130
rect 6391 1306 6425 1322
rect 6391 114 6425 130
rect 6569 1306 6603 1322
rect 6569 114 6603 130
rect 6747 1306 6781 1322
rect 6747 114 6781 130
rect 6925 1306 6959 1322
rect 6925 114 6959 130
rect 7103 1306 7137 1322
rect 7103 114 7137 130
rect 7281 1306 7315 1322
rect 7281 114 7315 130
rect 7459 1306 7493 1322
rect 7459 114 7493 130
rect 7637 1306 7671 1322
rect 7637 114 7671 130
rect 7815 1306 7849 1322
rect 7815 114 7849 130
rect 7993 1306 8027 1322
rect 7993 114 8027 130
rect -7981 37 -7965 71
rect -7877 37 -7861 71
rect -7803 37 -7787 71
rect -7699 37 -7683 71
rect -7625 37 -7609 71
rect -7521 37 -7505 71
rect -7447 37 -7431 71
rect -7343 37 -7327 71
rect -7269 37 -7253 71
rect -7165 37 -7149 71
rect -7091 37 -7075 71
rect -6987 37 -6971 71
rect -6913 37 -6897 71
rect -6809 37 -6793 71
rect -6735 37 -6719 71
rect -6631 37 -6615 71
rect -6557 37 -6541 71
rect -6453 37 -6437 71
rect -6379 37 -6363 71
rect -6275 37 -6259 71
rect -6201 37 -6185 71
rect -6097 37 -6081 71
rect -6023 37 -6007 71
rect -5919 37 -5903 71
rect -5845 37 -5829 71
rect -5741 37 -5725 71
rect -5667 37 -5651 71
rect -5563 37 -5547 71
rect -5489 37 -5473 71
rect -5385 37 -5369 71
rect -5311 37 -5295 71
rect -5207 37 -5191 71
rect -5133 37 -5117 71
rect -5029 37 -5013 71
rect -4955 37 -4939 71
rect -4851 37 -4835 71
rect -4777 37 -4761 71
rect -4673 37 -4657 71
rect -4599 37 -4583 71
rect -4495 37 -4479 71
rect -4421 37 -4405 71
rect -4317 37 -4301 71
rect -4243 37 -4227 71
rect -4139 37 -4123 71
rect -4065 37 -4049 71
rect -3961 37 -3945 71
rect -3887 37 -3871 71
rect -3783 37 -3767 71
rect -3709 37 -3693 71
rect -3605 37 -3589 71
rect -3531 37 -3515 71
rect -3427 37 -3411 71
rect -3353 37 -3337 71
rect -3249 37 -3233 71
rect -3175 37 -3159 71
rect -3071 37 -3055 71
rect -2997 37 -2981 71
rect -2893 37 -2877 71
rect -2819 37 -2803 71
rect -2715 37 -2699 71
rect -2641 37 -2625 71
rect -2537 37 -2521 71
rect -2463 37 -2447 71
rect -2359 37 -2343 71
rect -2285 37 -2269 71
rect -2181 37 -2165 71
rect -2107 37 -2091 71
rect -2003 37 -1987 71
rect -1929 37 -1913 71
rect -1825 37 -1809 71
rect -1751 37 -1735 71
rect -1647 37 -1631 71
rect -1573 37 -1557 71
rect -1469 37 -1453 71
rect -1395 37 -1379 71
rect -1291 37 -1275 71
rect -1217 37 -1201 71
rect -1113 37 -1097 71
rect -1039 37 -1023 71
rect -935 37 -919 71
rect -861 37 -845 71
rect -757 37 -741 71
rect -683 37 -667 71
rect -579 37 -563 71
rect -505 37 -489 71
rect -401 37 -385 71
rect -327 37 -311 71
rect -223 37 -207 71
rect -149 37 -133 71
rect -45 37 -29 71
rect 29 37 45 71
rect 133 37 149 71
rect 207 37 223 71
rect 311 37 327 71
rect 385 37 401 71
rect 489 37 505 71
rect 563 37 579 71
rect 667 37 683 71
rect 741 37 757 71
rect 845 37 861 71
rect 919 37 935 71
rect 1023 37 1039 71
rect 1097 37 1113 71
rect 1201 37 1217 71
rect 1275 37 1291 71
rect 1379 37 1395 71
rect 1453 37 1469 71
rect 1557 37 1573 71
rect 1631 37 1647 71
rect 1735 37 1751 71
rect 1809 37 1825 71
rect 1913 37 1929 71
rect 1987 37 2003 71
rect 2091 37 2107 71
rect 2165 37 2181 71
rect 2269 37 2285 71
rect 2343 37 2359 71
rect 2447 37 2463 71
rect 2521 37 2537 71
rect 2625 37 2641 71
rect 2699 37 2715 71
rect 2803 37 2819 71
rect 2877 37 2893 71
rect 2981 37 2997 71
rect 3055 37 3071 71
rect 3159 37 3175 71
rect 3233 37 3249 71
rect 3337 37 3353 71
rect 3411 37 3427 71
rect 3515 37 3531 71
rect 3589 37 3605 71
rect 3693 37 3709 71
rect 3767 37 3783 71
rect 3871 37 3887 71
rect 3945 37 3961 71
rect 4049 37 4065 71
rect 4123 37 4139 71
rect 4227 37 4243 71
rect 4301 37 4317 71
rect 4405 37 4421 71
rect 4479 37 4495 71
rect 4583 37 4599 71
rect 4657 37 4673 71
rect 4761 37 4777 71
rect 4835 37 4851 71
rect 4939 37 4955 71
rect 5013 37 5029 71
rect 5117 37 5133 71
rect 5191 37 5207 71
rect 5295 37 5311 71
rect 5369 37 5385 71
rect 5473 37 5489 71
rect 5547 37 5563 71
rect 5651 37 5667 71
rect 5725 37 5741 71
rect 5829 37 5845 71
rect 5903 37 5919 71
rect 6007 37 6023 71
rect 6081 37 6097 71
rect 6185 37 6201 71
rect 6259 37 6275 71
rect 6363 37 6379 71
rect 6437 37 6453 71
rect 6541 37 6557 71
rect 6615 37 6631 71
rect 6719 37 6735 71
rect 6793 37 6809 71
rect 6897 37 6913 71
rect 6971 37 6987 71
rect 7075 37 7091 71
rect 7149 37 7165 71
rect 7253 37 7269 71
rect 7327 37 7343 71
rect 7431 37 7447 71
rect 7505 37 7521 71
rect 7609 37 7625 71
rect 7683 37 7699 71
rect 7787 37 7803 71
rect 7861 37 7877 71
rect 7965 37 7981 71
rect -7981 -71 -7965 -37
rect -7877 -71 -7861 -37
rect -7803 -71 -7787 -37
rect -7699 -71 -7683 -37
rect -7625 -71 -7609 -37
rect -7521 -71 -7505 -37
rect -7447 -71 -7431 -37
rect -7343 -71 -7327 -37
rect -7269 -71 -7253 -37
rect -7165 -71 -7149 -37
rect -7091 -71 -7075 -37
rect -6987 -71 -6971 -37
rect -6913 -71 -6897 -37
rect -6809 -71 -6793 -37
rect -6735 -71 -6719 -37
rect -6631 -71 -6615 -37
rect -6557 -71 -6541 -37
rect -6453 -71 -6437 -37
rect -6379 -71 -6363 -37
rect -6275 -71 -6259 -37
rect -6201 -71 -6185 -37
rect -6097 -71 -6081 -37
rect -6023 -71 -6007 -37
rect -5919 -71 -5903 -37
rect -5845 -71 -5829 -37
rect -5741 -71 -5725 -37
rect -5667 -71 -5651 -37
rect -5563 -71 -5547 -37
rect -5489 -71 -5473 -37
rect -5385 -71 -5369 -37
rect -5311 -71 -5295 -37
rect -5207 -71 -5191 -37
rect -5133 -71 -5117 -37
rect -5029 -71 -5013 -37
rect -4955 -71 -4939 -37
rect -4851 -71 -4835 -37
rect -4777 -71 -4761 -37
rect -4673 -71 -4657 -37
rect -4599 -71 -4583 -37
rect -4495 -71 -4479 -37
rect -4421 -71 -4405 -37
rect -4317 -71 -4301 -37
rect -4243 -71 -4227 -37
rect -4139 -71 -4123 -37
rect -4065 -71 -4049 -37
rect -3961 -71 -3945 -37
rect -3887 -71 -3871 -37
rect -3783 -71 -3767 -37
rect -3709 -71 -3693 -37
rect -3605 -71 -3589 -37
rect -3531 -71 -3515 -37
rect -3427 -71 -3411 -37
rect -3353 -71 -3337 -37
rect -3249 -71 -3233 -37
rect -3175 -71 -3159 -37
rect -3071 -71 -3055 -37
rect -2997 -71 -2981 -37
rect -2893 -71 -2877 -37
rect -2819 -71 -2803 -37
rect -2715 -71 -2699 -37
rect -2641 -71 -2625 -37
rect -2537 -71 -2521 -37
rect -2463 -71 -2447 -37
rect -2359 -71 -2343 -37
rect -2285 -71 -2269 -37
rect -2181 -71 -2165 -37
rect -2107 -71 -2091 -37
rect -2003 -71 -1987 -37
rect -1929 -71 -1913 -37
rect -1825 -71 -1809 -37
rect -1751 -71 -1735 -37
rect -1647 -71 -1631 -37
rect -1573 -71 -1557 -37
rect -1469 -71 -1453 -37
rect -1395 -71 -1379 -37
rect -1291 -71 -1275 -37
rect -1217 -71 -1201 -37
rect -1113 -71 -1097 -37
rect -1039 -71 -1023 -37
rect -935 -71 -919 -37
rect -861 -71 -845 -37
rect -757 -71 -741 -37
rect -683 -71 -667 -37
rect -579 -71 -563 -37
rect -505 -71 -489 -37
rect -401 -71 -385 -37
rect -327 -71 -311 -37
rect -223 -71 -207 -37
rect -149 -71 -133 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 133 -71 149 -37
rect 207 -71 223 -37
rect 311 -71 327 -37
rect 385 -71 401 -37
rect 489 -71 505 -37
rect 563 -71 579 -37
rect 667 -71 683 -37
rect 741 -71 757 -37
rect 845 -71 861 -37
rect 919 -71 935 -37
rect 1023 -71 1039 -37
rect 1097 -71 1113 -37
rect 1201 -71 1217 -37
rect 1275 -71 1291 -37
rect 1379 -71 1395 -37
rect 1453 -71 1469 -37
rect 1557 -71 1573 -37
rect 1631 -71 1647 -37
rect 1735 -71 1751 -37
rect 1809 -71 1825 -37
rect 1913 -71 1929 -37
rect 1987 -71 2003 -37
rect 2091 -71 2107 -37
rect 2165 -71 2181 -37
rect 2269 -71 2285 -37
rect 2343 -71 2359 -37
rect 2447 -71 2463 -37
rect 2521 -71 2537 -37
rect 2625 -71 2641 -37
rect 2699 -71 2715 -37
rect 2803 -71 2819 -37
rect 2877 -71 2893 -37
rect 2981 -71 2997 -37
rect 3055 -71 3071 -37
rect 3159 -71 3175 -37
rect 3233 -71 3249 -37
rect 3337 -71 3353 -37
rect 3411 -71 3427 -37
rect 3515 -71 3531 -37
rect 3589 -71 3605 -37
rect 3693 -71 3709 -37
rect 3767 -71 3783 -37
rect 3871 -71 3887 -37
rect 3945 -71 3961 -37
rect 4049 -71 4065 -37
rect 4123 -71 4139 -37
rect 4227 -71 4243 -37
rect 4301 -71 4317 -37
rect 4405 -71 4421 -37
rect 4479 -71 4495 -37
rect 4583 -71 4599 -37
rect 4657 -71 4673 -37
rect 4761 -71 4777 -37
rect 4835 -71 4851 -37
rect 4939 -71 4955 -37
rect 5013 -71 5029 -37
rect 5117 -71 5133 -37
rect 5191 -71 5207 -37
rect 5295 -71 5311 -37
rect 5369 -71 5385 -37
rect 5473 -71 5489 -37
rect 5547 -71 5563 -37
rect 5651 -71 5667 -37
rect 5725 -71 5741 -37
rect 5829 -71 5845 -37
rect 5903 -71 5919 -37
rect 6007 -71 6023 -37
rect 6081 -71 6097 -37
rect 6185 -71 6201 -37
rect 6259 -71 6275 -37
rect 6363 -71 6379 -37
rect 6437 -71 6453 -37
rect 6541 -71 6557 -37
rect 6615 -71 6631 -37
rect 6719 -71 6735 -37
rect 6793 -71 6809 -37
rect 6897 -71 6913 -37
rect 6971 -71 6987 -37
rect 7075 -71 7091 -37
rect 7149 -71 7165 -37
rect 7253 -71 7269 -37
rect 7327 -71 7343 -37
rect 7431 -71 7447 -37
rect 7505 -71 7521 -37
rect 7609 -71 7625 -37
rect 7683 -71 7699 -37
rect 7787 -71 7803 -37
rect 7861 -71 7877 -37
rect 7965 -71 7981 -37
rect -8027 -130 -7993 -114
rect -8027 -1322 -7993 -1306
rect -7849 -130 -7815 -114
rect -7849 -1322 -7815 -1306
rect -7671 -130 -7637 -114
rect -7671 -1322 -7637 -1306
rect -7493 -130 -7459 -114
rect -7493 -1322 -7459 -1306
rect -7315 -130 -7281 -114
rect -7315 -1322 -7281 -1306
rect -7137 -130 -7103 -114
rect -7137 -1322 -7103 -1306
rect -6959 -130 -6925 -114
rect -6959 -1322 -6925 -1306
rect -6781 -130 -6747 -114
rect -6781 -1322 -6747 -1306
rect -6603 -130 -6569 -114
rect -6603 -1322 -6569 -1306
rect -6425 -130 -6391 -114
rect -6425 -1322 -6391 -1306
rect -6247 -130 -6213 -114
rect -6247 -1322 -6213 -1306
rect -6069 -130 -6035 -114
rect -6069 -1322 -6035 -1306
rect -5891 -130 -5857 -114
rect -5891 -1322 -5857 -1306
rect -5713 -130 -5679 -114
rect -5713 -1322 -5679 -1306
rect -5535 -130 -5501 -114
rect -5535 -1322 -5501 -1306
rect -5357 -130 -5323 -114
rect -5357 -1322 -5323 -1306
rect -5179 -130 -5145 -114
rect -5179 -1322 -5145 -1306
rect -5001 -130 -4967 -114
rect -5001 -1322 -4967 -1306
rect -4823 -130 -4789 -114
rect -4823 -1322 -4789 -1306
rect -4645 -130 -4611 -114
rect -4645 -1322 -4611 -1306
rect -4467 -130 -4433 -114
rect -4467 -1322 -4433 -1306
rect -4289 -130 -4255 -114
rect -4289 -1322 -4255 -1306
rect -4111 -130 -4077 -114
rect -4111 -1322 -4077 -1306
rect -3933 -130 -3899 -114
rect -3933 -1322 -3899 -1306
rect -3755 -130 -3721 -114
rect -3755 -1322 -3721 -1306
rect -3577 -130 -3543 -114
rect -3577 -1322 -3543 -1306
rect -3399 -130 -3365 -114
rect -3399 -1322 -3365 -1306
rect -3221 -130 -3187 -114
rect -3221 -1322 -3187 -1306
rect -3043 -130 -3009 -114
rect -3043 -1322 -3009 -1306
rect -2865 -130 -2831 -114
rect -2865 -1322 -2831 -1306
rect -2687 -130 -2653 -114
rect -2687 -1322 -2653 -1306
rect -2509 -130 -2475 -114
rect -2509 -1322 -2475 -1306
rect -2331 -130 -2297 -114
rect -2331 -1322 -2297 -1306
rect -2153 -130 -2119 -114
rect -2153 -1322 -2119 -1306
rect -1975 -130 -1941 -114
rect -1975 -1322 -1941 -1306
rect -1797 -130 -1763 -114
rect -1797 -1322 -1763 -1306
rect -1619 -130 -1585 -114
rect -1619 -1322 -1585 -1306
rect -1441 -130 -1407 -114
rect -1441 -1322 -1407 -1306
rect -1263 -130 -1229 -114
rect -1263 -1322 -1229 -1306
rect -1085 -130 -1051 -114
rect -1085 -1322 -1051 -1306
rect -907 -130 -873 -114
rect -907 -1322 -873 -1306
rect -729 -130 -695 -114
rect -729 -1322 -695 -1306
rect -551 -130 -517 -114
rect -551 -1322 -517 -1306
rect -373 -130 -339 -114
rect -373 -1322 -339 -1306
rect -195 -130 -161 -114
rect -195 -1322 -161 -1306
rect -17 -130 17 -114
rect -17 -1322 17 -1306
rect 161 -130 195 -114
rect 161 -1322 195 -1306
rect 339 -130 373 -114
rect 339 -1322 373 -1306
rect 517 -130 551 -114
rect 517 -1322 551 -1306
rect 695 -130 729 -114
rect 695 -1322 729 -1306
rect 873 -130 907 -114
rect 873 -1322 907 -1306
rect 1051 -130 1085 -114
rect 1051 -1322 1085 -1306
rect 1229 -130 1263 -114
rect 1229 -1322 1263 -1306
rect 1407 -130 1441 -114
rect 1407 -1322 1441 -1306
rect 1585 -130 1619 -114
rect 1585 -1322 1619 -1306
rect 1763 -130 1797 -114
rect 1763 -1322 1797 -1306
rect 1941 -130 1975 -114
rect 1941 -1322 1975 -1306
rect 2119 -130 2153 -114
rect 2119 -1322 2153 -1306
rect 2297 -130 2331 -114
rect 2297 -1322 2331 -1306
rect 2475 -130 2509 -114
rect 2475 -1322 2509 -1306
rect 2653 -130 2687 -114
rect 2653 -1322 2687 -1306
rect 2831 -130 2865 -114
rect 2831 -1322 2865 -1306
rect 3009 -130 3043 -114
rect 3009 -1322 3043 -1306
rect 3187 -130 3221 -114
rect 3187 -1322 3221 -1306
rect 3365 -130 3399 -114
rect 3365 -1322 3399 -1306
rect 3543 -130 3577 -114
rect 3543 -1322 3577 -1306
rect 3721 -130 3755 -114
rect 3721 -1322 3755 -1306
rect 3899 -130 3933 -114
rect 3899 -1322 3933 -1306
rect 4077 -130 4111 -114
rect 4077 -1322 4111 -1306
rect 4255 -130 4289 -114
rect 4255 -1322 4289 -1306
rect 4433 -130 4467 -114
rect 4433 -1322 4467 -1306
rect 4611 -130 4645 -114
rect 4611 -1322 4645 -1306
rect 4789 -130 4823 -114
rect 4789 -1322 4823 -1306
rect 4967 -130 5001 -114
rect 4967 -1322 5001 -1306
rect 5145 -130 5179 -114
rect 5145 -1322 5179 -1306
rect 5323 -130 5357 -114
rect 5323 -1322 5357 -1306
rect 5501 -130 5535 -114
rect 5501 -1322 5535 -1306
rect 5679 -130 5713 -114
rect 5679 -1322 5713 -1306
rect 5857 -130 5891 -114
rect 5857 -1322 5891 -1306
rect 6035 -130 6069 -114
rect 6035 -1322 6069 -1306
rect 6213 -130 6247 -114
rect 6213 -1322 6247 -1306
rect 6391 -130 6425 -114
rect 6391 -1322 6425 -1306
rect 6569 -130 6603 -114
rect 6569 -1322 6603 -1306
rect 6747 -130 6781 -114
rect 6747 -1322 6781 -1306
rect 6925 -130 6959 -114
rect 6925 -1322 6959 -1306
rect 7103 -130 7137 -114
rect 7103 -1322 7137 -1306
rect 7281 -130 7315 -114
rect 7281 -1322 7315 -1306
rect 7459 -130 7493 -114
rect 7459 -1322 7493 -1306
rect 7637 -130 7671 -114
rect 7637 -1322 7671 -1306
rect 7815 -130 7849 -114
rect 7815 -1322 7849 -1306
rect 7993 -130 8027 -114
rect 7993 -1322 8027 -1306
rect -7981 -1399 -7965 -1365
rect -7877 -1399 -7861 -1365
rect -7803 -1399 -7787 -1365
rect -7699 -1399 -7683 -1365
rect -7625 -1399 -7609 -1365
rect -7521 -1399 -7505 -1365
rect -7447 -1399 -7431 -1365
rect -7343 -1399 -7327 -1365
rect -7269 -1399 -7253 -1365
rect -7165 -1399 -7149 -1365
rect -7091 -1399 -7075 -1365
rect -6987 -1399 -6971 -1365
rect -6913 -1399 -6897 -1365
rect -6809 -1399 -6793 -1365
rect -6735 -1399 -6719 -1365
rect -6631 -1399 -6615 -1365
rect -6557 -1399 -6541 -1365
rect -6453 -1399 -6437 -1365
rect -6379 -1399 -6363 -1365
rect -6275 -1399 -6259 -1365
rect -6201 -1399 -6185 -1365
rect -6097 -1399 -6081 -1365
rect -6023 -1399 -6007 -1365
rect -5919 -1399 -5903 -1365
rect -5845 -1399 -5829 -1365
rect -5741 -1399 -5725 -1365
rect -5667 -1399 -5651 -1365
rect -5563 -1399 -5547 -1365
rect -5489 -1399 -5473 -1365
rect -5385 -1399 -5369 -1365
rect -5311 -1399 -5295 -1365
rect -5207 -1399 -5191 -1365
rect -5133 -1399 -5117 -1365
rect -5029 -1399 -5013 -1365
rect -4955 -1399 -4939 -1365
rect -4851 -1399 -4835 -1365
rect -4777 -1399 -4761 -1365
rect -4673 -1399 -4657 -1365
rect -4599 -1399 -4583 -1365
rect -4495 -1399 -4479 -1365
rect -4421 -1399 -4405 -1365
rect -4317 -1399 -4301 -1365
rect -4243 -1399 -4227 -1365
rect -4139 -1399 -4123 -1365
rect -4065 -1399 -4049 -1365
rect -3961 -1399 -3945 -1365
rect -3887 -1399 -3871 -1365
rect -3783 -1399 -3767 -1365
rect -3709 -1399 -3693 -1365
rect -3605 -1399 -3589 -1365
rect -3531 -1399 -3515 -1365
rect -3427 -1399 -3411 -1365
rect -3353 -1399 -3337 -1365
rect -3249 -1399 -3233 -1365
rect -3175 -1399 -3159 -1365
rect -3071 -1399 -3055 -1365
rect -2997 -1399 -2981 -1365
rect -2893 -1399 -2877 -1365
rect -2819 -1399 -2803 -1365
rect -2715 -1399 -2699 -1365
rect -2641 -1399 -2625 -1365
rect -2537 -1399 -2521 -1365
rect -2463 -1399 -2447 -1365
rect -2359 -1399 -2343 -1365
rect -2285 -1399 -2269 -1365
rect -2181 -1399 -2165 -1365
rect -2107 -1399 -2091 -1365
rect -2003 -1399 -1987 -1365
rect -1929 -1399 -1913 -1365
rect -1825 -1399 -1809 -1365
rect -1751 -1399 -1735 -1365
rect -1647 -1399 -1631 -1365
rect -1573 -1399 -1557 -1365
rect -1469 -1399 -1453 -1365
rect -1395 -1399 -1379 -1365
rect -1291 -1399 -1275 -1365
rect -1217 -1399 -1201 -1365
rect -1113 -1399 -1097 -1365
rect -1039 -1399 -1023 -1365
rect -935 -1399 -919 -1365
rect -861 -1399 -845 -1365
rect -757 -1399 -741 -1365
rect -683 -1399 -667 -1365
rect -579 -1399 -563 -1365
rect -505 -1399 -489 -1365
rect -401 -1399 -385 -1365
rect -327 -1399 -311 -1365
rect -223 -1399 -207 -1365
rect -149 -1399 -133 -1365
rect -45 -1399 -29 -1365
rect 29 -1399 45 -1365
rect 133 -1399 149 -1365
rect 207 -1399 223 -1365
rect 311 -1399 327 -1365
rect 385 -1399 401 -1365
rect 489 -1399 505 -1365
rect 563 -1399 579 -1365
rect 667 -1399 683 -1365
rect 741 -1399 757 -1365
rect 845 -1399 861 -1365
rect 919 -1399 935 -1365
rect 1023 -1399 1039 -1365
rect 1097 -1399 1113 -1365
rect 1201 -1399 1217 -1365
rect 1275 -1399 1291 -1365
rect 1379 -1399 1395 -1365
rect 1453 -1399 1469 -1365
rect 1557 -1399 1573 -1365
rect 1631 -1399 1647 -1365
rect 1735 -1399 1751 -1365
rect 1809 -1399 1825 -1365
rect 1913 -1399 1929 -1365
rect 1987 -1399 2003 -1365
rect 2091 -1399 2107 -1365
rect 2165 -1399 2181 -1365
rect 2269 -1399 2285 -1365
rect 2343 -1399 2359 -1365
rect 2447 -1399 2463 -1365
rect 2521 -1399 2537 -1365
rect 2625 -1399 2641 -1365
rect 2699 -1399 2715 -1365
rect 2803 -1399 2819 -1365
rect 2877 -1399 2893 -1365
rect 2981 -1399 2997 -1365
rect 3055 -1399 3071 -1365
rect 3159 -1399 3175 -1365
rect 3233 -1399 3249 -1365
rect 3337 -1399 3353 -1365
rect 3411 -1399 3427 -1365
rect 3515 -1399 3531 -1365
rect 3589 -1399 3605 -1365
rect 3693 -1399 3709 -1365
rect 3767 -1399 3783 -1365
rect 3871 -1399 3887 -1365
rect 3945 -1399 3961 -1365
rect 4049 -1399 4065 -1365
rect 4123 -1399 4139 -1365
rect 4227 -1399 4243 -1365
rect 4301 -1399 4317 -1365
rect 4405 -1399 4421 -1365
rect 4479 -1399 4495 -1365
rect 4583 -1399 4599 -1365
rect 4657 -1399 4673 -1365
rect 4761 -1399 4777 -1365
rect 4835 -1399 4851 -1365
rect 4939 -1399 4955 -1365
rect 5013 -1399 5029 -1365
rect 5117 -1399 5133 -1365
rect 5191 -1399 5207 -1365
rect 5295 -1399 5311 -1365
rect 5369 -1399 5385 -1365
rect 5473 -1399 5489 -1365
rect 5547 -1399 5563 -1365
rect 5651 -1399 5667 -1365
rect 5725 -1399 5741 -1365
rect 5829 -1399 5845 -1365
rect 5903 -1399 5919 -1365
rect 6007 -1399 6023 -1365
rect 6081 -1399 6097 -1365
rect 6185 -1399 6201 -1365
rect 6259 -1399 6275 -1365
rect 6363 -1399 6379 -1365
rect 6437 -1399 6453 -1365
rect 6541 -1399 6557 -1365
rect 6615 -1399 6631 -1365
rect 6719 -1399 6735 -1365
rect 6793 -1399 6809 -1365
rect 6897 -1399 6913 -1365
rect 6971 -1399 6987 -1365
rect 7075 -1399 7091 -1365
rect 7149 -1399 7165 -1365
rect 7253 -1399 7269 -1365
rect 7327 -1399 7343 -1365
rect 7431 -1399 7447 -1365
rect 7505 -1399 7521 -1365
rect 7609 -1399 7625 -1365
rect 7683 -1399 7699 -1365
rect 7787 -1399 7803 -1365
rect 7861 -1399 7877 -1365
rect 7965 -1399 7981 -1365
rect -8141 -1467 -8107 -1405
rect 8107 -1467 8141 -1405
rect -8141 -1501 -8045 -1467
rect 8045 -1501 8141 -1467
<< viali >>
rect -7965 1365 -7877 1399
rect -7787 1365 -7699 1399
rect -7609 1365 -7521 1399
rect -7431 1365 -7343 1399
rect -7253 1365 -7165 1399
rect -7075 1365 -6987 1399
rect -6897 1365 -6809 1399
rect -6719 1365 -6631 1399
rect -6541 1365 -6453 1399
rect -6363 1365 -6275 1399
rect -6185 1365 -6097 1399
rect -6007 1365 -5919 1399
rect -5829 1365 -5741 1399
rect -5651 1365 -5563 1399
rect -5473 1365 -5385 1399
rect -5295 1365 -5207 1399
rect -5117 1365 -5029 1399
rect -4939 1365 -4851 1399
rect -4761 1365 -4673 1399
rect -4583 1365 -4495 1399
rect -4405 1365 -4317 1399
rect -4227 1365 -4139 1399
rect -4049 1365 -3961 1399
rect -3871 1365 -3783 1399
rect -3693 1365 -3605 1399
rect -3515 1365 -3427 1399
rect -3337 1365 -3249 1399
rect -3159 1365 -3071 1399
rect -2981 1365 -2893 1399
rect -2803 1365 -2715 1399
rect -2625 1365 -2537 1399
rect -2447 1365 -2359 1399
rect -2269 1365 -2181 1399
rect -2091 1365 -2003 1399
rect -1913 1365 -1825 1399
rect -1735 1365 -1647 1399
rect -1557 1365 -1469 1399
rect -1379 1365 -1291 1399
rect -1201 1365 -1113 1399
rect -1023 1365 -935 1399
rect -845 1365 -757 1399
rect -667 1365 -579 1399
rect -489 1365 -401 1399
rect -311 1365 -223 1399
rect -133 1365 -45 1399
rect 45 1365 133 1399
rect 223 1365 311 1399
rect 401 1365 489 1399
rect 579 1365 667 1399
rect 757 1365 845 1399
rect 935 1365 1023 1399
rect 1113 1365 1201 1399
rect 1291 1365 1379 1399
rect 1469 1365 1557 1399
rect 1647 1365 1735 1399
rect 1825 1365 1913 1399
rect 2003 1365 2091 1399
rect 2181 1365 2269 1399
rect 2359 1365 2447 1399
rect 2537 1365 2625 1399
rect 2715 1365 2803 1399
rect 2893 1365 2981 1399
rect 3071 1365 3159 1399
rect 3249 1365 3337 1399
rect 3427 1365 3515 1399
rect 3605 1365 3693 1399
rect 3783 1365 3871 1399
rect 3961 1365 4049 1399
rect 4139 1365 4227 1399
rect 4317 1365 4405 1399
rect 4495 1365 4583 1399
rect 4673 1365 4761 1399
rect 4851 1365 4939 1399
rect 5029 1365 5117 1399
rect 5207 1365 5295 1399
rect 5385 1365 5473 1399
rect 5563 1365 5651 1399
rect 5741 1365 5829 1399
rect 5919 1365 6007 1399
rect 6097 1365 6185 1399
rect 6275 1365 6363 1399
rect 6453 1365 6541 1399
rect 6631 1365 6719 1399
rect 6809 1365 6897 1399
rect 6987 1365 7075 1399
rect 7165 1365 7253 1399
rect 7343 1365 7431 1399
rect 7521 1365 7609 1399
rect 7699 1365 7787 1399
rect 7877 1365 7965 1399
rect -8027 130 -7993 1306
rect -7849 130 -7815 1306
rect -7671 130 -7637 1306
rect -7493 130 -7459 1306
rect -7315 130 -7281 1306
rect -7137 130 -7103 1306
rect -6959 130 -6925 1306
rect -6781 130 -6747 1306
rect -6603 130 -6569 1306
rect -6425 130 -6391 1306
rect -6247 130 -6213 1306
rect -6069 130 -6035 1306
rect -5891 130 -5857 1306
rect -5713 130 -5679 1306
rect -5535 130 -5501 1306
rect -5357 130 -5323 1306
rect -5179 130 -5145 1306
rect -5001 130 -4967 1306
rect -4823 130 -4789 1306
rect -4645 130 -4611 1306
rect -4467 130 -4433 1306
rect -4289 130 -4255 1306
rect -4111 130 -4077 1306
rect -3933 130 -3899 1306
rect -3755 130 -3721 1306
rect -3577 130 -3543 1306
rect -3399 130 -3365 1306
rect -3221 130 -3187 1306
rect -3043 130 -3009 1306
rect -2865 130 -2831 1306
rect -2687 130 -2653 1306
rect -2509 130 -2475 1306
rect -2331 130 -2297 1306
rect -2153 130 -2119 1306
rect -1975 130 -1941 1306
rect -1797 130 -1763 1306
rect -1619 130 -1585 1306
rect -1441 130 -1407 1306
rect -1263 130 -1229 1306
rect -1085 130 -1051 1306
rect -907 130 -873 1306
rect -729 130 -695 1306
rect -551 130 -517 1306
rect -373 130 -339 1306
rect -195 130 -161 1306
rect -17 130 17 1306
rect 161 130 195 1306
rect 339 130 373 1306
rect 517 130 551 1306
rect 695 130 729 1306
rect 873 130 907 1306
rect 1051 130 1085 1306
rect 1229 130 1263 1306
rect 1407 130 1441 1306
rect 1585 130 1619 1306
rect 1763 130 1797 1306
rect 1941 130 1975 1306
rect 2119 130 2153 1306
rect 2297 130 2331 1306
rect 2475 130 2509 1306
rect 2653 130 2687 1306
rect 2831 130 2865 1306
rect 3009 130 3043 1306
rect 3187 130 3221 1306
rect 3365 130 3399 1306
rect 3543 130 3577 1306
rect 3721 130 3755 1306
rect 3899 130 3933 1306
rect 4077 130 4111 1306
rect 4255 130 4289 1306
rect 4433 130 4467 1306
rect 4611 130 4645 1306
rect 4789 130 4823 1306
rect 4967 130 5001 1306
rect 5145 130 5179 1306
rect 5323 130 5357 1306
rect 5501 130 5535 1306
rect 5679 130 5713 1306
rect 5857 130 5891 1306
rect 6035 130 6069 1306
rect 6213 130 6247 1306
rect 6391 130 6425 1306
rect 6569 130 6603 1306
rect 6747 130 6781 1306
rect 6925 130 6959 1306
rect 7103 130 7137 1306
rect 7281 130 7315 1306
rect 7459 130 7493 1306
rect 7637 130 7671 1306
rect 7815 130 7849 1306
rect 7993 130 8027 1306
rect -7965 37 -7877 71
rect -7787 37 -7699 71
rect -7609 37 -7521 71
rect -7431 37 -7343 71
rect -7253 37 -7165 71
rect -7075 37 -6987 71
rect -6897 37 -6809 71
rect -6719 37 -6631 71
rect -6541 37 -6453 71
rect -6363 37 -6275 71
rect -6185 37 -6097 71
rect -6007 37 -5919 71
rect -5829 37 -5741 71
rect -5651 37 -5563 71
rect -5473 37 -5385 71
rect -5295 37 -5207 71
rect -5117 37 -5029 71
rect -4939 37 -4851 71
rect -4761 37 -4673 71
rect -4583 37 -4495 71
rect -4405 37 -4317 71
rect -4227 37 -4139 71
rect -4049 37 -3961 71
rect -3871 37 -3783 71
rect -3693 37 -3605 71
rect -3515 37 -3427 71
rect -3337 37 -3249 71
rect -3159 37 -3071 71
rect -2981 37 -2893 71
rect -2803 37 -2715 71
rect -2625 37 -2537 71
rect -2447 37 -2359 71
rect -2269 37 -2181 71
rect -2091 37 -2003 71
rect -1913 37 -1825 71
rect -1735 37 -1647 71
rect -1557 37 -1469 71
rect -1379 37 -1291 71
rect -1201 37 -1113 71
rect -1023 37 -935 71
rect -845 37 -757 71
rect -667 37 -579 71
rect -489 37 -401 71
rect -311 37 -223 71
rect -133 37 -45 71
rect 45 37 133 71
rect 223 37 311 71
rect 401 37 489 71
rect 579 37 667 71
rect 757 37 845 71
rect 935 37 1023 71
rect 1113 37 1201 71
rect 1291 37 1379 71
rect 1469 37 1557 71
rect 1647 37 1735 71
rect 1825 37 1913 71
rect 2003 37 2091 71
rect 2181 37 2269 71
rect 2359 37 2447 71
rect 2537 37 2625 71
rect 2715 37 2803 71
rect 2893 37 2981 71
rect 3071 37 3159 71
rect 3249 37 3337 71
rect 3427 37 3515 71
rect 3605 37 3693 71
rect 3783 37 3871 71
rect 3961 37 4049 71
rect 4139 37 4227 71
rect 4317 37 4405 71
rect 4495 37 4583 71
rect 4673 37 4761 71
rect 4851 37 4939 71
rect 5029 37 5117 71
rect 5207 37 5295 71
rect 5385 37 5473 71
rect 5563 37 5651 71
rect 5741 37 5829 71
rect 5919 37 6007 71
rect 6097 37 6185 71
rect 6275 37 6363 71
rect 6453 37 6541 71
rect 6631 37 6719 71
rect 6809 37 6897 71
rect 6987 37 7075 71
rect 7165 37 7253 71
rect 7343 37 7431 71
rect 7521 37 7609 71
rect 7699 37 7787 71
rect 7877 37 7965 71
rect -7965 -71 -7877 -37
rect -7787 -71 -7699 -37
rect -7609 -71 -7521 -37
rect -7431 -71 -7343 -37
rect -7253 -71 -7165 -37
rect -7075 -71 -6987 -37
rect -6897 -71 -6809 -37
rect -6719 -71 -6631 -37
rect -6541 -71 -6453 -37
rect -6363 -71 -6275 -37
rect -6185 -71 -6097 -37
rect -6007 -71 -5919 -37
rect -5829 -71 -5741 -37
rect -5651 -71 -5563 -37
rect -5473 -71 -5385 -37
rect -5295 -71 -5207 -37
rect -5117 -71 -5029 -37
rect -4939 -71 -4851 -37
rect -4761 -71 -4673 -37
rect -4583 -71 -4495 -37
rect -4405 -71 -4317 -37
rect -4227 -71 -4139 -37
rect -4049 -71 -3961 -37
rect -3871 -71 -3783 -37
rect -3693 -71 -3605 -37
rect -3515 -71 -3427 -37
rect -3337 -71 -3249 -37
rect -3159 -71 -3071 -37
rect -2981 -71 -2893 -37
rect -2803 -71 -2715 -37
rect -2625 -71 -2537 -37
rect -2447 -71 -2359 -37
rect -2269 -71 -2181 -37
rect -2091 -71 -2003 -37
rect -1913 -71 -1825 -37
rect -1735 -71 -1647 -37
rect -1557 -71 -1469 -37
rect -1379 -71 -1291 -37
rect -1201 -71 -1113 -37
rect -1023 -71 -935 -37
rect -845 -71 -757 -37
rect -667 -71 -579 -37
rect -489 -71 -401 -37
rect -311 -71 -223 -37
rect -133 -71 -45 -37
rect 45 -71 133 -37
rect 223 -71 311 -37
rect 401 -71 489 -37
rect 579 -71 667 -37
rect 757 -71 845 -37
rect 935 -71 1023 -37
rect 1113 -71 1201 -37
rect 1291 -71 1379 -37
rect 1469 -71 1557 -37
rect 1647 -71 1735 -37
rect 1825 -71 1913 -37
rect 2003 -71 2091 -37
rect 2181 -71 2269 -37
rect 2359 -71 2447 -37
rect 2537 -71 2625 -37
rect 2715 -71 2803 -37
rect 2893 -71 2981 -37
rect 3071 -71 3159 -37
rect 3249 -71 3337 -37
rect 3427 -71 3515 -37
rect 3605 -71 3693 -37
rect 3783 -71 3871 -37
rect 3961 -71 4049 -37
rect 4139 -71 4227 -37
rect 4317 -71 4405 -37
rect 4495 -71 4583 -37
rect 4673 -71 4761 -37
rect 4851 -71 4939 -37
rect 5029 -71 5117 -37
rect 5207 -71 5295 -37
rect 5385 -71 5473 -37
rect 5563 -71 5651 -37
rect 5741 -71 5829 -37
rect 5919 -71 6007 -37
rect 6097 -71 6185 -37
rect 6275 -71 6363 -37
rect 6453 -71 6541 -37
rect 6631 -71 6719 -37
rect 6809 -71 6897 -37
rect 6987 -71 7075 -37
rect 7165 -71 7253 -37
rect 7343 -71 7431 -37
rect 7521 -71 7609 -37
rect 7699 -71 7787 -37
rect 7877 -71 7965 -37
rect -8027 -1306 -7993 -130
rect -7849 -1306 -7815 -130
rect -7671 -1306 -7637 -130
rect -7493 -1306 -7459 -130
rect -7315 -1306 -7281 -130
rect -7137 -1306 -7103 -130
rect -6959 -1306 -6925 -130
rect -6781 -1306 -6747 -130
rect -6603 -1306 -6569 -130
rect -6425 -1306 -6391 -130
rect -6247 -1306 -6213 -130
rect -6069 -1306 -6035 -130
rect -5891 -1306 -5857 -130
rect -5713 -1306 -5679 -130
rect -5535 -1306 -5501 -130
rect -5357 -1306 -5323 -130
rect -5179 -1306 -5145 -130
rect -5001 -1306 -4967 -130
rect -4823 -1306 -4789 -130
rect -4645 -1306 -4611 -130
rect -4467 -1306 -4433 -130
rect -4289 -1306 -4255 -130
rect -4111 -1306 -4077 -130
rect -3933 -1306 -3899 -130
rect -3755 -1306 -3721 -130
rect -3577 -1306 -3543 -130
rect -3399 -1306 -3365 -130
rect -3221 -1306 -3187 -130
rect -3043 -1306 -3009 -130
rect -2865 -1306 -2831 -130
rect -2687 -1306 -2653 -130
rect -2509 -1306 -2475 -130
rect -2331 -1306 -2297 -130
rect -2153 -1306 -2119 -130
rect -1975 -1306 -1941 -130
rect -1797 -1306 -1763 -130
rect -1619 -1306 -1585 -130
rect -1441 -1306 -1407 -130
rect -1263 -1306 -1229 -130
rect -1085 -1306 -1051 -130
rect -907 -1306 -873 -130
rect -729 -1306 -695 -130
rect -551 -1306 -517 -130
rect -373 -1306 -339 -130
rect -195 -1306 -161 -130
rect -17 -1306 17 -130
rect 161 -1306 195 -130
rect 339 -1306 373 -130
rect 517 -1306 551 -130
rect 695 -1306 729 -130
rect 873 -1306 907 -130
rect 1051 -1306 1085 -130
rect 1229 -1306 1263 -130
rect 1407 -1306 1441 -130
rect 1585 -1306 1619 -130
rect 1763 -1306 1797 -130
rect 1941 -1306 1975 -130
rect 2119 -1306 2153 -130
rect 2297 -1306 2331 -130
rect 2475 -1306 2509 -130
rect 2653 -1306 2687 -130
rect 2831 -1306 2865 -130
rect 3009 -1306 3043 -130
rect 3187 -1306 3221 -130
rect 3365 -1306 3399 -130
rect 3543 -1306 3577 -130
rect 3721 -1306 3755 -130
rect 3899 -1306 3933 -130
rect 4077 -1306 4111 -130
rect 4255 -1306 4289 -130
rect 4433 -1306 4467 -130
rect 4611 -1306 4645 -130
rect 4789 -1306 4823 -130
rect 4967 -1306 5001 -130
rect 5145 -1306 5179 -130
rect 5323 -1306 5357 -130
rect 5501 -1306 5535 -130
rect 5679 -1306 5713 -130
rect 5857 -1306 5891 -130
rect 6035 -1306 6069 -130
rect 6213 -1306 6247 -130
rect 6391 -1306 6425 -130
rect 6569 -1306 6603 -130
rect 6747 -1306 6781 -130
rect 6925 -1306 6959 -130
rect 7103 -1306 7137 -130
rect 7281 -1306 7315 -130
rect 7459 -1306 7493 -130
rect 7637 -1306 7671 -130
rect 7815 -1306 7849 -130
rect 7993 -1306 8027 -130
rect -7965 -1399 -7877 -1365
rect -7787 -1399 -7699 -1365
rect -7609 -1399 -7521 -1365
rect -7431 -1399 -7343 -1365
rect -7253 -1399 -7165 -1365
rect -7075 -1399 -6987 -1365
rect -6897 -1399 -6809 -1365
rect -6719 -1399 -6631 -1365
rect -6541 -1399 -6453 -1365
rect -6363 -1399 -6275 -1365
rect -6185 -1399 -6097 -1365
rect -6007 -1399 -5919 -1365
rect -5829 -1399 -5741 -1365
rect -5651 -1399 -5563 -1365
rect -5473 -1399 -5385 -1365
rect -5295 -1399 -5207 -1365
rect -5117 -1399 -5029 -1365
rect -4939 -1399 -4851 -1365
rect -4761 -1399 -4673 -1365
rect -4583 -1399 -4495 -1365
rect -4405 -1399 -4317 -1365
rect -4227 -1399 -4139 -1365
rect -4049 -1399 -3961 -1365
rect -3871 -1399 -3783 -1365
rect -3693 -1399 -3605 -1365
rect -3515 -1399 -3427 -1365
rect -3337 -1399 -3249 -1365
rect -3159 -1399 -3071 -1365
rect -2981 -1399 -2893 -1365
rect -2803 -1399 -2715 -1365
rect -2625 -1399 -2537 -1365
rect -2447 -1399 -2359 -1365
rect -2269 -1399 -2181 -1365
rect -2091 -1399 -2003 -1365
rect -1913 -1399 -1825 -1365
rect -1735 -1399 -1647 -1365
rect -1557 -1399 -1469 -1365
rect -1379 -1399 -1291 -1365
rect -1201 -1399 -1113 -1365
rect -1023 -1399 -935 -1365
rect -845 -1399 -757 -1365
rect -667 -1399 -579 -1365
rect -489 -1399 -401 -1365
rect -311 -1399 -223 -1365
rect -133 -1399 -45 -1365
rect 45 -1399 133 -1365
rect 223 -1399 311 -1365
rect 401 -1399 489 -1365
rect 579 -1399 667 -1365
rect 757 -1399 845 -1365
rect 935 -1399 1023 -1365
rect 1113 -1399 1201 -1365
rect 1291 -1399 1379 -1365
rect 1469 -1399 1557 -1365
rect 1647 -1399 1735 -1365
rect 1825 -1399 1913 -1365
rect 2003 -1399 2091 -1365
rect 2181 -1399 2269 -1365
rect 2359 -1399 2447 -1365
rect 2537 -1399 2625 -1365
rect 2715 -1399 2803 -1365
rect 2893 -1399 2981 -1365
rect 3071 -1399 3159 -1365
rect 3249 -1399 3337 -1365
rect 3427 -1399 3515 -1365
rect 3605 -1399 3693 -1365
rect 3783 -1399 3871 -1365
rect 3961 -1399 4049 -1365
rect 4139 -1399 4227 -1365
rect 4317 -1399 4405 -1365
rect 4495 -1399 4583 -1365
rect 4673 -1399 4761 -1365
rect 4851 -1399 4939 -1365
rect 5029 -1399 5117 -1365
rect 5207 -1399 5295 -1365
rect 5385 -1399 5473 -1365
rect 5563 -1399 5651 -1365
rect 5741 -1399 5829 -1365
rect 5919 -1399 6007 -1365
rect 6097 -1399 6185 -1365
rect 6275 -1399 6363 -1365
rect 6453 -1399 6541 -1365
rect 6631 -1399 6719 -1365
rect 6809 -1399 6897 -1365
rect 6987 -1399 7075 -1365
rect 7165 -1399 7253 -1365
rect 7343 -1399 7431 -1365
rect 7521 -1399 7609 -1365
rect 7699 -1399 7787 -1365
rect 7877 -1399 7965 -1365
<< metal1 >>
rect -7977 1399 -7865 1405
rect -7977 1365 -7965 1399
rect -7877 1365 -7865 1399
rect -7977 1359 -7865 1365
rect -7799 1399 -7687 1405
rect -7799 1365 -7787 1399
rect -7699 1365 -7687 1399
rect -7799 1359 -7687 1365
rect -7621 1399 -7509 1405
rect -7621 1365 -7609 1399
rect -7521 1365 -7509 1399
rect -7621 1359 -7509 1365
rect -7443 1399 -7331 1405
rect -7443 1365 -7431 1399
rect -7343 1365 -7331 1399
rect -7443 1359 -7331 1365
rect -7265 1399 -7153 1405
rect -7265 1365 -7253 1399
rect -7165 1365 -7153 1399
rect -7265 1359 -7153 1365
rect -7087 1399 -6975 1405
rect -7087 1365 -7075 1399
rect -6987 1365 -6975 1399
rect -7087 1359 -6975 1365
rect -6909 1399 -6797 1405
rect -6909 1365 -6897 1399
rect -6809 1365 -6797 1399
rect -6909 1359 -6797 1365
rect -6731 1399 -6619 1405
rect -6731 1365 -6719 1399
rect -6631 1365 -6619 1399
rect -6731 1359 -6619 1365
rect -6553 1399 -6441 1405
rect -6553 1365 -6541 1399
rect -6453 1365 -6441 1399
rect -6553 1359 -6441 1365
rect -6375 1399 -6263 1405
rect -6375 1365 -6363 1399
rect -6275 1365 -6263 1399
rect -6375 1359 -6263 1365
rect -6197 1399 -6085 1405
rect -6197 1365 -6185 1399
rect -6097 1365 -6085 1399
rect -6197 1359 -6085 1365
rect -6019 1399 -5907 1405
rect -6019 1365 -6007 1399
rect -5919 1365 -5907 1399
rect -6019 1359 -5907 1365
rect -5841 1399 -5729 1405
rect -5841 1365 -5829 1399
rect -5741 1365 -5729 1399
rect -5841 1359 -5729 1365
rect -5663 1399 -5551 1405
rect -5663 1365 -5651 1399
rect -5563 1365 -5551 1399
rect -5663 1359 -5551 1365
rect -5485 1399 -5373 1405
rect -5485 1365 -5473 1399
rect -5385 1365 -5373 1399
rect -5485 1359 -5373 1365
rect -5307 1399 -5195 1405
rect -5307 1365 -5295 1399
rect -5207 1365 -5195 1399
rect -5307 1359 -5195 1365
rect -5129 1399 -5017 1405
rect -5129 1365 -5117 1399
rect -5029 1365 -5017 1399
rect -5129 1359 -5017 1365
rect -4951 1399 -4839 1405
rect -4951 1365 -4939 1399
rect -4851 1365 -4839 1399
rect -4951 1359 -4839 1365
rect -4773 1399 -4661 1405
rect -4773 1365 -4761 1399
rect -4673 1365 -4661 1399
rect -4773 1359 -4661 1365
rect -4595 1399 -4483 1405
rect -4595 1365 -4583 1399
rect -4495 1365 -4483 1399
rect -4595 1359 -4483 1365
rect -4417 1399 -4305 1405
rect -4417 1365 -4405 1399
rect -4317 1365 -4305 1399
rect -4417 1359 -4305 1365
rect -4239 1399 -4127 1405
rect -4239 1365 -4227 1399
rect -4139 1365 -4127 1399
rect -4239 1359 -4127 1365
rect -4061 1399 -3949 1405
rect -4061 1365 -4049 1399
rect -3961 1365 -3949 1399
rect -4061 1359 -3949 1365
rect -3883 1399 -3771 1405
rect -3883 1365 -3871 1399
rect -3783 1365 -3771 1399
rect -3883 1359 -3771 1365
rect -3705 1399 -3593 1405
rect -3705 1365 -3693 1399
rect -3605 1365 -3593 1399
rect -3705 1359 -3593 1365
rect -3527 1399 -3415 1405
rect -3527 1365 -3515 1399
rect -3427 1365 -3415 1399
rect -3527 1359 -3415 1365
rect -3349 1399 -3237 1405
rect -3349 1365 -3337 1399
rect -3249 1365 -3237 1399
rect -3349 1359 -3237 1365
rect -3171 1399 -3059 1405
rect -3171 1365 -3159 1399
rect -3071 1365 -3059 1399
rect -3171 1359 -3059 1365
rect -2993 1399 -2881 1405
rect -2993 1365 -2981 1399
rect -2893 1365 -2881 1399
rect -2993 1359 -2881 1365
rect -2815 1399 -2703 1405
rect -2815 1365 -2803 1399
rect -2715 1365 -2703 1399
rect -2815 1359 -2703 1365
rect -2637 1399 -2525 1405
rect -2637 1365 -2625 1399
rect -2537 1365 -2525 1399
rect -2637 1359 -2525 1365
rect -2459 1399 -2347 1405
rect -2459 1365 -2447 1399
rect -2359 1365 -2347 1399
rect -2459 1359 -2347 1365
rect -2281 1399 -2169 1405
rect -2281 1365 -2269 1399
rect -2181 1365 -2169 1399
rect -2281 1359 -2169 1365
rect -2103 1399 -1991 1405
rect -2103 1365 -2091 1399
rect -2003 1365 -1991 1399
rect -2103 1359 -1991 1365
rect -1925 1399 -1813 1405
rect -1925 1365 -1913 1399
rect -1825 1365 -1813 1399
rect -1925 1359 -1813 1365
rect -1747 1399 -1635 1405
rect -1747 1365 -1735 1399
rect -1647 1365 -1635 1399
rect -1747 1359 -1635 1365
rect -1569 1399 -1457 1405
rect -1569 1365 -1557 1399
rect -1469 1365 -1457 1399
rect -1569 1359 -1457 1365
rect -1391 1399 -1279 1405
rect -1391 1365 -1379 1399
rect -1291 1365 -1279 1399
rect -1391 1359 -1279 1365
rect -1213 1399 -1101 1405
rect -1213 1365 -1201 1399
rect -1113 1365 -1101 1399
rect -1213 1359 -1101 1365
rect -1035 1399 -923 1405
rect -1035 1365 -1023 1399
rect -935 1365 -923 1399
rect -1035 1359 -923 1365
rect -857 1399 -745 1405
rect -857 1365 -845 1399
rect -757 1365 -745 1399
rect -857 1359 -745 1365
rect -679 1399 -567 1405
rect -679 1365 -667 1399
rect -579 1365 -567 1399
rect -679 1359 -567 1365
rect -501 1399 -389 1405
rect -501 1365 -489 1399
rect -401 1365 -389 1399
rect -501 1359 -389 1365
rect -323 1399 -211 1405
rect -323 1365 -311 1399
rect -223 1365 -211 1399
rect -323 1359 -211 1365
rect -145 1399 -33 1405
rect -145 1365 -133 1399
rect -45 1365 -33 1399
rect -145 1359 -33 1365
rect 33 1399 145 1405
rect 33 1365 45 1399
rect 133 1365 145 1399
rect 33 1359 145 1365
rect 211 1399 323 1405
rect 211 1365 223 1399
rect 311 1365 323 1399
rect 211 1359 323 1365
rect 389 1399 501 1405
rect 389 1365 401 1399
rect 489 1365 501 1399
rect 389 1359 501 1365
rect 567 1399 679 1405
rect 567 1365 579 1399
rect 667 1365 679 1399
rect 567 1359 679 1365
rect 745 1399 857 1405
rect 745 1365 757 1399
rect 845 1365 857 1399
rect 745 1359 857 1365
rect 923 1399 1035 1405
rect 923 1365 935 1399
rect 1023 1365 1035 1399
rect 923 1359 1035 1365
rect 1101 1399 1213 1405
rect 1101 1365 1113 1399
rect 1201 1365 1213 1399
rect 1101 1359 1213 1365
rect 1279 1399 1391 1405
rect 1279 1365 1291 1399
rect 1379 1365 1391 1399
rect 1279 1359 1391 1365
rect 1457 1399 1569 1405
rect 1457 1365 1469 1399
rect 1557 1365 1569 1399
rect 1457 1359 1569 1365
rect 1635 1399 1747 1405
rect 1635 1365 1647 1399
rect 1735 1365 1747 1399
rect 1635 1359 1747 1365
rect 1813 1399 1925 1405
rect 1813 1365 1825 1399
rect 1913 1365 1925 1399
rect 1813 1359 1925 1365
rect 1991 1399 2103 1405
rect 1991 1365 2003 1399
rect 2091 1365 2103 1399
rect 1991 1359 2103 1365
rect 2169 1399 2281 1405
rect 2169 1365 2181 1399
rect 2269 1365 2281 1399
rect 2169 1359 2281 1365
rect 2347 1399 2459 1405
rect 2347 1365 2359 1399
rect 2447 1365 2459 1399
rect 2347 1359 2459 1365
rect 2525 1399 2637 1405
rect 2525 1365 2537 1399
rect 2625 1365 2637 1399
rect 2525 1359 2637 1365
rect 2703 1399 2815 1405
rect 2703 1365 2715 1399
rect 2803 1365 2815 1399
rect 2703 1359 2815 1365
rect 2881 1399 2993 1405
rect 2881 1365 2893 1399
rect 2981 1365 2993 1399
rect 2881 1359 2993 1365
rect 3059 1399 3171 1405
rect 3059 1365 3071 1399
rect 3159 1365 3171 1399
rect 3059 1359 3171 1365
rect 3237 1399 3349 1405
rect 3237 1365 3249 1399
rect 3337 1365 3349 1399
rect 3237 1359 3349 1365
rect 3415 1399 3527 1405
rect 3415 1365 3427 1399
rect 3515 1365 3527 1399
rect 3415 1359 3527 1365
rect 3593 1399 3705 1405
rect 3593 1365 3605 1399
rect 3693 1365 3705 1399
rect 3593 1359 3705 1365
rect 3771 1399 3883 1405
rect 3771 1365 3783 1399
rect 3871 1365 3883 1399
rect 3771 1359 3883 1365
rect 3949 1399 4061 1405
rect 3949 1365 3961 1399
rect 4049 1365 4061 1399
rect 3949 1359 4061 1365
rect 4127 1399 4239 1405
rect 4127 1365 4139 1399
rect 4227 1365 4239 1399
rect 4127 1359 4239 1365
rect 4305 1399 4417 1405
rect 4305 1365 4317 1399
rect 4405 1365 4417 1399
rect 4305 1359 4417 1365
rect 4483 1399 4595 1405
rect 4483 1365 4495 1399
rect 4583 1365 4595 1399
rect 4483 1359 4595 1365
rect 4661 1399 4773 1405
rect 4661 1365 4673 1399
rect 4761 1365 4773 1399
rect 4661 1359 4773 1365
rect 4839 1399 4951 1405
rect 4839 1365 4851 1399
rect 4939 1365 4951 1399
rect 4839 1359 4951 1365
rect 5017 1399 5129 1405
rect 5017 1365 5029 1399
rect 5117 1365 5129 1399
rect 5017 1359 5129 1365
rect 5195 1399 5307 1405
rect 5195 1365 5207 1399
rect 5295 1365 5307 1399
rect 5195 1359 5307 1365
rect 5373 1399 5485 1405
rect 5373 1365 5385 1399
rect 5473 1365 5485 1399
rect 5373 1359 5485 1365
rect 5551 1399 5663 1405
rect 5551 1365 5563 1399
rect 5651 1365 5663 1399
rect 5551 1359 5663 1365
rect 5729 1399 5841 1405
rect 5729 1365 5741 1399
rect 5829 1365 5841 1399
rect 5729 1359 5841 1365
rect 5907 1399 6019 1405
rect 5907 1365 5919 1399
rect 6007 1365 6019 1399
rect 5907 1359 6019 1365
rect 6085 1399 6197 1405
rect 6085 1365 6097 1399
rect 6185 1365 6197 1399
rect 6085 1359 6197 1365
rect 6263 1399 6375 1405
rect 6263 1365 6275 1399
rect 6363 1365 6375 1399
rect 6263 1359 6375 1365
rect 6441 1399 6553 1405
rect 6441 1365 6453 1399
rect 6541 1365 6553 1399
rect 6441 1359 6553 1365
rect 6619 1399 6731 1405
rect 6619 1365 6631 1399
rect 6719 1365 6731 1399
rect 6619 1359 6731 1365
rect 6797 1399 6909 1405
rect 6797 1365 6809 1399
rect 6897 1365 6909 1399
rect 6797 1359 6909 1365
rect 6975 1399 7087 1405
rect 6975 1365 6987 1399
rect 7075 1365 7087 1399
rect 6975 1359 7087 1365
rect 7153 1399 7265 1405
rect 7153 1365 7165 1399
rect 7253 1365 7265 1399
rect 7153 1359 7265 1365
rect 7331 1399 7443 1405
rect 7331 1365 7343 1399
rect 7431 1365 7443 1399
rect 7331 1359 7443 1365
rect 7509 1399 7621 1405
rect 7509 1365 7521 1399
rect 7609 1365 7621 1399
rect 7509 1359 7621 1365
rect 7687 1399 7799 1405
rect 7687 1365 7699 1399
rect 7787 1365 7799 1399
rect 7687 1359 7799 1365
rect 7865 1399 7977 1405
rect 7865 1365 7877 1399
rect 7965 1365 7977 1399
rect 7865 1359 7977 1365
rect -8033 1306 -7987 1318
rect -8033 130 -8027 1306
rect -7993 130 -7987 1306
rect -8033 118 -7987 130
rect -7855 1306 -7809 1318
rect -7855 130 -7849 1306
rect -7815 130 -7809 1306
rect -7855 118 -7809 130
rect -7677 1306 -7631 1318
rect -7677 130 -7671 1306
rect -7637 130 -7631 1306
rect -7677 118 -7631 130
rect -7499 1306 -7453 1318
rect -7499 130 -7493 1306
rect -7459 130 -7453 1306
rect -7499 118 -7453 130
rect -7321 1306 -7275 1318
rect -7321 130 -7315 1306
rect -7281 130 -7275 1306
rect -7321 118 -7275 130
rect -7143 1306 -7097 1318
rect -7143 130 -7137 1306
rect -7103 130 -7097 1306
rect -7143 118 -7097 130
rect -6965 1306 -6919 1318
rect -6965 130 -6959 1306
rect -6925 130 -6919 1306
rect -6965 118 -6919 130
rect -6787 1306 -6741 1318
rect -6787 130 -6781 1306
rect -6747 130 -6741 1306
rect -6787 118 -6741 130
rect -6609 1306 -6563 1318
rect -6609 130 -6603 1306
rect -6569 130 -6563 1306
rect -6609 118 -6563 130
rect -6431 1306 -6385 1318
rect -6431 130 -6425 1306
rect -6391 130 -6385 1306
rect -6431 118 -6385 130
rect -6253 1306 -6207 1318
rect -6253 130 -6247 1306
rect -6213 130 -6207 1306
rect -6253 118 -6207 130
rect -6075 1306 -6029 1318
rect -6075 130 -6069 1306
rect -6035 130 -6029 1306
rect -6075 118 -6029 130
rect -5897 1306 -5851 1318
rect -5897 130 -5891 1306
rect -5857 130 -5851 1306
rect -5897 118 -5851 130
rect -5719 1306 -5673 1318
rect -5719 130 -5713 1306
rect -5679 130 -5673 1306
rect -5719 118 -5673 130
rect -5541 1306 -5495 1318
rect -5541 130 -5535 1306
rect -5501 130 -5495 1306
rect -5541 118 -5495 130
rect -5363 1306 -5317 1318
rect -5363 130 -5357 1306
rect -5323 130 -5317 1306
rect -5363 118 -5317 130
rect -5185 1306 -5139 1318
rect -5185 130 -5179 1306
rect -5145 130 -5139 1306
rect -5185 118 -5139 130
rect -5007 1306 -4961 1318
rect -5007 130 -5001 1306
rect -4967 130 -4961 1306
rect -5007 118 -4961 130
rect -4829 1306 -4783 1318
rect -4829 130 -4823 1306
rect -4789 130 -4783 1306
rect -4829 118 -4783 130
rect -4651 1306 -4605 1318
rect -4651 130 -4645 1306
rect -4611 130 -4605 1306
rect -4651 118 -4605 130
rect -4473 1306 -4427 1318
rect -4473 130 -4467 1306
rect -4433 130 -4427 1306
rect -4473 118 -4427 130
rect -4295 1306 -4249 1318
rect -4295 130 -4289 1306
rect -4255 130 -4249 1306
rect -4295 118 -4249 130
rect -4117 1306 -4071 1318
rect -4117 130 -4111 1306
rect -4077 130 -4071 1306
rect -4117 118 -4071 130
rect -3939 1306 -3893 1318
rect -3939 130 -3933 1306
rect -3899 130 -3893 1306
rect -3939 118 -3893 130
rect -3761 1306 -3715 1318
rect -3761 130 -3755 1306
rect -3721 130 -3715 1306
rect -3761 118 -3715 130
rect -3583 1306 -3537 1318
rect -3583 130 -3577 1306
rect -3543 130 -3537 1306
rect -3583 118 -3537 130
rect -3405 1306 -3359 1318
rect -3405 130 -3399 1306
rect -3365 130 -3359 1306
rect -3405 118 -3359 130
rect -3227 1306 -3181 1318
rect -3227 130 -3221 1306
rect -3187 130 -3181 1306
rect -3227 118 -3181 130
rect -3049 1306 -3003 1318
rect -3049 130 -3043 1306
rect -3009 130 -3003 1306
rect -3049 118 -3003 130
rect -2871 1306 -2825 1318
rect -2871 130 -2865 1306
rect -2831 130 -2825 1306
rect -2871 118 -2825 130
rect -2693 1306 -2647 1318
rect -2693 130 -2687 1306
rect -2653 130 -2647 1306
rect -2693 118 -2647 130
rect -2515 1306 -2469 1318
rect -2515 130 -2509 1306
rect -2475 130 -2469 1306
rect -2515 118 -2469 130
rect -2337 1306 -2291 1318
rect -2337 130 -2331 1306
rect -2297 130 -2291 1306
rect -2337 118 -2291 130
rect -2159 1306 -2113 1318
rect -2159 130 -2153 1306
rect -2119 130 -2113 1306
rect -2159 118 -2113 130
rect -1981 1306 -1935 1318
rect -1981 130 -1975 1306
rect -1941 130 -1935 1306
rect -1981 118 -1935 130
rect -1803 1306 -1757 1318
rect -1803 130 -1797 1306
rect -1763 130 -1757 1306
rect -1803 118 -1757 130
rect -1625 1306 -1579 1318
rect -1625 130 -1619 1306
rect -1585 130 -1579 1306
rect -1625 118 -1579 130
rect -1447 1306 -1401 1318
rect -1447 130 -1441 1306
rect -1407 130 -1401 1306
rect -1447 118 -1401 130
rect -1269 1306 -1223 1318
rect -1269 130 -1263 1306
rect -1229 130 -1223 1306
rect -1269 118 -1223 130
rect -1091 1306 -1045 1318
rect -1091 130 -1085 1306
rect -1051 130 -1045 1306
rect -1091 118 -1045 130
rect -913 1306 -867 1318
rect -913 130 -907 1306
rect -873 130 -867 1306
rect -913 118 -867 130
rect -735 1306 -689 1318
rect -735 130 -729 1306
rect -695 130 -689 1306
rect -735 118 -689 130
rect -557 1306 -511 1318
rect -557 130 -551 1306
rect -517 130 -511 1306
rect -557 118 -511 130
rect -379 1306 -333 1318
rect -379 130 -373 1306
rect -339 130 -333 1306
rect -379 118 -333 130
rect -201 1306 -155 1318
rect -201 130 -195 1306
rect -161 130 -155 1306
rect -201 118 -155 130
rect -23 1306 23 1318
rect -23 130 -17 1306
rect 17 130 23 1306
rect -23 118 23 130
rect 155 1306 201 1318
rect 155 130 161 1306
rect 195 130 201 1306
rect 155 118 201 130
rect 333 1306 379 1318
rect 333 130 339 1306
rect 373 130 379 1306
rect 333 118 379 130
rect 511 1306 557 1318
rect 511 130 517 1306
rect 551 130 557 1306
rect 511 118 557 130
rect 689 1306 735 1318
rect 689 130 695 1306
rect 729 130 735 1306
rect 689 118 735 130
rect 867 1306 913 1318
rect 867 130 873 1306
rect 907 130 913 1306
rect 867 118 913 130
rect 1045 1306 1091 1318
rect 1045 130 1051 1306
rect 1085 130 1091 1306
rect 1045 118 1091 130
rect 1223 1306 1269 1318
rect 1223 130 1229 1306
rect 1263 130 1269 1306
rect 1223 118 1269 130
rect 1401 1306 1447 1318
rect 1401 130 1407 1306
rect 1441 130 1447 1306
rect 1401 118 1447 130
rect 1579 1306 1625 1318
rect 1579 130 1585 1306
rect 1619 130 1625 1306
rect 1579 118 1625 130
rect 1757 1306 1803 1318
rect 1757 130 1763 1306
rect 1797 130 1803 1306
rect 1757 118 1803 130
rect 1935 1306 1981 1318
rect 1935 130 1941 1306
rect 1975 130 1981 1306
rect 1935 118 1981 130
rect 2113 1306 2159 1318
rect 2113 130 2119 1306
rect 2153 130 2159 1306
rect 2113 118 2159 130
rect 2291 1306 2337 1318
rect 2291 130 2297 1306
rect 2331 130 2337 1306
rect 2291 118 2337 130
rect 2469 1306 2515 1318
rect 2469 130 2475 1306
rect 2509 130 2515 1306
rect 2469 118 2515 130
rect 2647 1306 2693 1318
rect 2647 130 2653 1306
rect 2687 130 2693 1306
rect 2647 118 2693 130
rect 2825 1306 2871 1318
rect 2825 130 2831 1306
rect 2865 130 2871 1306
rect 2825 118 2871 130
rect 3003 1306 3049 1318
rect 3003 130 3009 1306
rect 3043 130 3049 1306
rect 3003 118 3049 130
rect 3181 1306 3227 1318
rect 3181 130 3187 1306
rect 3221 130 3227 1306
rect 3181 118 3227 130
rect 3359 1306 3405 1318
rect 3359 130 3365 1306
rect 3399 130 3405 1306
rect 3359 118 3405 130
rect 3537 1306 3583 1318
rect 3537 130 3543 1306
rect 3577 130 3583 1306
rect 3537 118 3583 130
rect 3715 1306 3761 1318
rect 3715 130 3721 1306
rect 3755 130 3761 1306
rect 3715 118 3761 130
rect 3893 1306 3939 1318
rect 3893 130 3899 1306
rect 3933 130 3939 1306
rect 3893 118 3939 130
rect 4071 1306 4117 1318
rect 4071 130 4077 1306
rect 4111 130 4117 1306
rect 4071 118 4117 130
rect 4249 1306 4295 1318
rect 4249 130 4255 1306
rect 4289 130 4295 1306
rect 4249 118 4295 130
rect 4427 1306 4473 1318
rect 4427 130 4433 1306
rect 4467 130 4473 1306
rect 4427 118 4473 130
rect 4605 1306 4651 1318
rect 4605 130 4611 1306
rect 4645 130 4651 1306
rect 4605 118 4651 130
rect 4783 1306 4829 1318
rect 4783 130 4789 1306
rect 4823 130 4829 1306
rect 4783 118 4829 130
rect 4961 1306 5007 1318
rect 4961 130 4967 1306
rect 5001 130 5007 1306
rect 4961 118 5007 130
rect 5139 1306 5185 1318
rect 5139 130 5145 1306
rect 5179 130 5185 1306
rect 5139 118 5185 130
rect 5317 1306 5363 1318
rect 5317 130 5323 1306
rect 5357 130 5363 1306
rect 5317 118 5363 130
rect 5495 1306 5541 1318
rect 5495 130 5501 1306
rect 5535 130 5541 1306
rect 5495 118 5541 130
rect 5673 1306 5719 1318
rect 5673 130 5679 1306
rect 5713 130 5719 1306
rect 5673 118 5719 130
rect 5851 1306 5897 1318
rect 5851 130 5857 1306
rect 5891 130 5897 1306
rect 5851 118 5897 130
rect 6029 1306 6075 1318
rect 6029 130 6035 1306
rect 6069 130 6075 1306
rect 6029 118 6075 130
rect 6207 1306 6253 1318
rect 6207 130 6213 1306
rect 6247 130 6253 1306
rect 6207 118 6253 130
rect 6385 1306 6431 1318
rect 6385 130 6391 1306
rect 6425 130 6431 1306
rect 6385 118 6431 130
rect 6563 1306 6609 1318
rect 6563 130 6569 1306
rect 6603 130 6609 1306
rect 6563 118 6609 130
rect 6741 1306 6787 1318
rect 6741 130 6747 1306
rect 6781 130 6787 1306
rect 6741 118 6787 130
rect 6919 1306 6965 1318
rect 6919 130 6925 1306
rect 6959 130 6965 1306
rect 6919 118 6965 130
rect 7097 1306 7143 1318
rect 7097 130 7103 1306
rect 7137 130 7143 1306
rect 7097 118 7143 130
rect 7275 1306 7321 1318
rect 7275 130 7281 1306
rect 7315 130 7321 1306
rect 7275 118 7321 130
rect 7453 1306 7499 1318
rect 7453 130 7459 1306
rect 7493 130 7499 1306
rect 7453 118 7499 130
rect 7631 1306 7677 1318
rect 7631 130 7637 1306
rect 7671 130 7677 1306
rect 7631 118 7677 130
rect 7809 1306 7855 1318
rect 7809 130 7815 1306
rect 7849 130 7855 1306
rect 7809 118 7855 130
rect 7987 1306 8033 1318
rect 7987 130 7993 1306
rect 8027 130 8033 1306
rect 7987 118 8033 130
rect -7977 71 -7865 77
rect -7977 37 -7965 71
rect -7877 37 -7865 71
rect -7977 31 -7865 37
rect -7799 71 -7687 77
rect -7799 37 -7787 71
rect -7699 37 -7687 71
rect -7799 31 -7687 37
rect -7621 71 -7509 77
rect -7621 37 -7609 71
rect -7521 37 -7509 71
rect -7621 31 -7509 37
rect -7443 71 -7331 77
rect -7443 37 -7431 71
rect -7343 37 -7331 71
rect -7443 31 -7331 37
rect -7265 71 -7153 77
rect -7265 37 -7253 71
rect -7165 37 -7153 71
rect -7265 31 -7153 37
rect -7087 71 -6975 77
rect -7087 37 -7075 71
rect -6987 37 -6975 71
rect -7087 31 -6975 37
rect -6909 71 -6797 77
rect -6909 37 -6897 71
rect -6809 37 -6797 71
rect -6909 31 -6797 37
rect -6731 71 -6619 77
rect -6731 37 -6719 71
rect -6631 37 -6619 71
rect -6731 31 -6619 37
rect -6553 71 -6441 77
rect -6553 37 -6541 71
rect -6453 37 -6441 71
rect -6553 31 -6441 37
rect -6375 71 -6263 77
rect -6375 37 -6363 71
rect -6275 37 -6263 71
rect -6375 31 -6263 37
rect -6197 71 -6085 77
rect -6197 37 -6185 71
rect -6097 37 -6085 71
rect -6197 31 -6085 37
rect -6019 71 -5907 77
rect -6019 37 -6007 71
rect -5919 37 -5907 71
rect -6019 31 -5907 37
rect -5841 71 -5729 77
rect -5841 37 -5829 71
rect -5741 37 -5729 71
rect -5841 31 -5729 37
rect -5663 71 -5551 77
rect -5663 37 -5651 71
rect -5563 37 -5551 71
rect -5663 31 -5551 37
rect -5485 71 -5373 77
rect -5485 37 -5473 71
rect -5385 37 -5373 71
rect -5485 31 -5373 37
rect -5307 71 -5195 77
rect -5307 37 -5295 71
rect -5207 37 -5195 71
rect -5307 31 -5195 37
rect -5129 71 -5017 77
rect -5129 37 -5117 71
rect -5029 37 -5017 71
rect -5129 31 -5017 37
rect -4951 71 -4839 77
rect -4951 37 -4939 71
rect -4851 37 -4839 71
rect -4951 31 -4839 37
rect -4773 71 -4661 77
rect -4773 37 -4761 71
rect -4673 37 -4661 71
rect -4773 31 -4661 37
rect -4595 71 -4483 77
rect -4595 37 -4583 71
rect -4495 37 -4483 71
rect -4595 31 -4483 37
rect -4417 71 -4305 77
rect -4417 37 -4405 71
rect -4317 37 -4305 71
rect -4417 31 -4305 37
rect -4239 71 -4127 77
rect -4239 37 -4227 71
rect -4139 37 -4127 71
rect -4239 31 -4127 37
rect -4061 71 -3949 77
rect -4061 37 -4049 71
rect -3961 37 -3949 71
rect -4061 31 -3949 37
rect -3883 71 -3771 77
rect -3883 37 -3871 71
rect -3783 37 -3771 71
rect -3883 31 -3771 37
rect -3705 71 -3593 77
rect -3705 37 -3693 71
rect -3605 37 -3593 71
rect -3705 31 -3593 37
rect -3527 71 -3415 77
rect -3527 37 -3515 71
rect -3427 37 -3415 71
rect -3527 31 -3415 37
rect -3349 71 -3237 77
rect -3349 37 -3337 71
rect -3249 37 -3237 71
rect -3349 31 -3237 37
rect -3171 71 -3059 77
rect -3171 37 -3159 71
rect -3071 37 -3059 71
rect -3171 31 -3059 37
rect -2993 71 -2881 77
rect -2993 37 -2981 71
rect -2893 37 -2881 71
rect -2993 31 -2881 37
rect -2815 71 -2703 77
rect -2815 37 -2803 71
rect -2715 37 -2703 71
rect -2815 31 -2703 37
rect -2637 71 -2525 77
rect -2637 37 -2625 71
rect -2537 37 -2525 71
rect -2637 31 -2525 37
rect -2459 71 -2347 77
rect -2459 37 -2447 71
rect -2359 37 -2347 71
rect -2459 31 -2347 37
rect -2281 71 -2169 77
rect -2281 37 -2269 71
rect -2181 37 -2169 71
rect -2281 31 -2169 37
rect -2103 71 -1991 77
rect -2103 37 -2091 71
rect -2003 37 -1991 71
rect -2103 31 -1991 37
rect -1925 71 -1813 77
rect -1925 37 -1913 71
rect -1825 37 -1813 71
rect -1925 31 -1813 37
rect -1747 71 -1635 77
rect -1747 37 -1735 71
rect -1647 37 -1635 71
rect -1747 31 -1635 37
rect -1569 71 -1457 77
rect -1569 37 -1557 71
rect -1469 37 -1457 71
rect -1569 31 -1457 37
rect -1391 71 -1279 77
rect -1391 37 -1379 71
rect -1291 37 -1279 71
rect -1391 31 -1279 37
rect -1213 71 -1101 77
rect -1213 37 -1201 71
rect -1113 37 -1101 71
rect -1213 31 -1101 37
rect -1035 71 -923 77
rect -1035 37 -1023 71
rect -935 37 -923 71
rect -1035 31 -923 37
rect -857 71 -745 77
rect -857 37 -845 71
rect -757 37 -745 71
rect -857 31 -745 37
rect -679 71 -567 77
rect -679 37 -667 71
rect -579 37 -567 71
rect -679 31 -567 37
rect -501 71 -389 77
rect -501 37 -489 71
rect -401 37 -389 71
rect -501 31 -389 37
rect -323 71 -211 77
rect -323 37 -311 71
rect -223 37 -211 71
rect -323 31 -211 37
rect -145 71 -33 77
rect -145 37 -133 71
rect -45 37 -33 71
rect -145 31 -33 37
rect 33 71 145 77
rect 33 37 45 71
rect 133 37 145 71
rect 33 31 145 37
rect 211 71 323 77
rect 211 37 223 71
rect 311 37 323 71
rect 211 31 323 37
rect 389 71 501 77
rect 389 37 401 71
rect 489 37 501 71
rect 389 31 501 37
rect 567 71 679 77
rect 567 37 579 71
rect 667 37 679 71
rect 567 31 679 37
rect 745 71 857 77
rect 745 37 757 71
rect 845 37 857 71
rect 745 31 857 37
rect 923 71 1035 77
rect 923 37 935 71
rect 1023 37 1035 71
rect 923 31 1035 37
rect 1101 71 1213 77
rect 1101 37 1113 71
rect 1201 37 1213 71
rect 1101 31 1213 37
rect 1279 71 1391 77
rect 1279 37 1291 71
rect 1379 37 1391 71
rect 1279 31 1391 37
rect 1457 71 1569 77
rect 1457 37 1469 71
rect 1557 37 1569 71
rect 1457 31 1569 37
rect 1635 71 1747 77
rect 1635 37 1647 71
rect 1735 37 1747 71
rect 1635 31 1747 37
rect 1813 71 1925 77
rect 1813 37 1825 71
rect 1913 37 1925 71
rect 1813 31 1925 37
rect 1991 71 2103 77
rect 1991 37 2003 71
rect 2091 37 2103 71
rect 1991 31 2103 37
rect 2169 71 2281 77
rect 2169 37 2181 71
rect 2269 37 2281 71
rect 2169 31 2281 37
rect 2347 71 2459 77
rect 2347 37 2359 71
rect 2447 37 2459 71
rect 2347 31 2459 37
rect 2525 71 2637 77
rect 2525 37 2537 71
rect 2625 37 2637 71
rect 2525 31 2637 37
rect 2703 71 2815 77
rect 2703 37 2715 71
rect 2803 37 2815 71
rect 2703 31 2815 37
rect 2881 71 2993 77
rect 2881 37 2893 71
rect 2981 37 2993 71
rect 2881 31 2993 37
rect 3059 71 3171 77
rect 3059 37 3071 71
rect 3159 37 3171 71
rect 3059 31 3171 37
rect 3237 71 3349 77
rect 3237 37 3249 71
rect 3337 37 3349 71
rect 3237 31 3349 37
rect 3415 71 3527 77
rect 3415 37 3427 71
rect 3515 37 3527 71
rect 3415 31 3527 37
rect 3593 71 3705 77
rect 3593 37 3605 71
rect 3693 37 3705 71
rect 3593 31 3705 37
rect 3771 71 3883 77
rect 3771 37 3783 71
rect 3871 37 3883 71
rect 3771 31 3883 37
rect 3949 71 4061 77
rect 3949 37 3961 71
rect 4049 37 4061 71
rect 3949 31 4061 37
rect 4127 71 4239 77
rect 4127 37 4139 71
rect 4227 37 4239 71
rect 4127 31 4239 37
rect 4305 71 4417 77
rect 4305 37 4317 71
rect 4405 37 4417 71
rect 4305 31 4417 37
rect 4483 71 4595 77
rect 4483 37 4495 71
rect 4583 37 4595 71
rect 4483 31 4595 37
rect 4661 71 4773 77
rect 4661 37 4673 71
rect 4761 37 4773 71
rect 4661 31 4773 37
rect 4839 71 4951 77
rect 4839 37 4851 71
rect 4939 37 4951 71
rect 4839 31 4951 37
rect 5017 71 5129 77
rect 5017 37 5029 71
rect 5117 37 5129 71
rect 5017 31 5129 37
rect 5195 71 5307 77
rect 5195 37 5207 71
rect 5295 37 5307 71
rect 5195 31 5307 37
rect 5373 71 5485 77
rect 5373 37 5385 71
rect 5473 37 5485 71
rect 5373 31 5485 37
rect 5551 71 5663 77
rect 5551 37 5563 71
rect 5651 37 5663 71
rect 5551 31 5663 37
rect 5729 71 5841 77
rect 5729 37 5741 71
rect 5829 37 5841 71
rect 5729 31 5841 37
rect 5907 71 6019 77
rect 5907 37 5919 71
rect 6007 37 6019 71
rect 5907 31 6019 37
rect 6085 71 6197 77
rect 6085 37 6097 71
rect 6185 37 6197 71
rect 6085 31 6197 37
rect 6263 71 6375 77
rect 6263 37 6275 71
rect 6363 37 6375 71
rect 6263 31 6375 37
rect 6441 71 6553 77
rect 6441 37 6453 71
rect 6541 37 6553 71
rect 6441 31 6553 37
rect 6619 71 6731 77
rect 6619 37 6631 71
rect 6719 37 6731 71
rect 6619 31 6731 37
rect 6797 71 6909 77
rect 6797 37 6809 71
rect 6897 37 6909 71
rect 6797 31 6909 37
rect 6975 71 7087 77
rect 6975 37 6987 71
rect 7075 37 7087 71
rect 6975 31 7087 37
rect 7153 71 7265 77
rect 7153 37 7165 71
rect 7253 37 7265 71
rect 7153 31 7265 37
rect 7331 71 7443 77
rect 7331 37 7343 71
rect 7431 37 7443 71
rect 7331 31 7443 37
rect 7509 71 7621 77
rect 7509 37 7521 71
rect 7609 37 7621 71
rect 7509 31 7621 37
rect 7687 71 7799 77
rect 7687 37 7699 71
rect 7787 37 7799 71
rect 7687 31 7799 37
rect 7865 71 7977 77
rect 7865 37 7877 71
rect 7965 37 7977 71
rect 7865 31 7977 37
rect -7977 -37 -7865 -31
rect -7977 -71 -7965 -37
rect -7877 -71 -7865 -37
rect -7977 -77 -7865 -71
rect -7799 -37 -7687 -31
rect -7799 -71 -7787 -37
rect -7699 -71 -7687 -37
rect -7799 -77 -7687 -71
rect -7621 -37 -7509 -31
rect -7621 -71 -7609 -37
rect -7521 -71 -7509 -37
rect -7621 -77 -7509 -71
rect -7443 -37 -7331 -31
rect -7443 -71 -7431 -37
rect -7343 -71 -7331 -37
rect -7443 -77 -7331 -71
rect -7265 -37 -7153 -31
rect -7265 -71 -7253 -37
rect -7165 -71 -7153 -37
rect -7265 -77 -7153 -71
rect -7087 -37 -6975 -31
rect -7087 -71 -7075 -37
rect -6987 -71 -6975 -37
rect -7087 -77 -6975 -71
rect -6909 -37 -6797 -31
rect -6909 -71 -6897 -37
rect -6809 -71 -6797 -37
rect -6909 -77 -6797 -71
rect -6731 -37 -6619 -31
rect -6731 -71 -6719 -37
rect -6631 -71 -6619 -37
rect -6731 -77 -6619 -71
rect -6553 -37 -6441 -31
rect -6553 -71 -6541 -37
rect -6453 -71 -6441 -37
rect -6553 -77 -6441 -71
rect -6375 -37 -6263 -31
rect -6375 -71 -6363 -37
rect -6275 -71 -6263 -37
rect -6375 -77 -6263 -71
rect -6197 -37 -6085 -31
rect -6197 -71 -6185 -37
rect -6097 -71 -6085 -37
rect -6197 -77 -6085 -71
rect -6019 -37 -5907 -31
rect -6019 -71 -6007 -37
rect -5919 -71 -5907 -37
rect -6019 -77 -5907 -71
rect -5841 -37 -5729 -31
rect -5841 -71 -5829 -37
rect -5741 -71 -5729 -37
rect -5841 -77 -5729 -71
rect -5663 -37 -5551 -31
rect -5663 -71 -5651 -37
rect -5563 -71 -5551 -37
rect -5663 -77 -5551 -71
rect -5485 -37 -5373 -31
rect -5485 -71 -5473 -37
rect -5385 -71 -5373 -37
rect -5485 -77 -5373 -71
rect -5307 -37 -5195 -31
rect -5307 -71 -5295 -37
rect -5207 -71 -5195 -37
rect -5307 -77 -5195 -71
rect -5129 -37 -5017 -31
rect -5129 -71 -5117 -37
rect -5029 -71 -5017 -37
rect -5129 -77 -5017 -71
rect -4951 -37 -4839 -31
rect -4951 -71 -4939 -37
rect -4851 -71 -4839 -37
rect -4951 -77 -4839 -71
rect -4773 -37 -4661 -31
rect -4773 -71 -4761 -37
rect -4673 -71 -4661 -37
rect -4773 -77 -4661 -71
rect -4595 -37 -4483 -31
rect -4595 -71 -4583 -37
rect -4495 -71 -4483 -37
rect -4595 -77 -4483 -71
rect -4417 -37 -4305 -31
rect -4417 -71 -4405 -37
rect -4317 -71 -4305 -37
rect -4417 -77 -4305 -71
rect -4239 -37 -4127 -31
rect -4239 -71 -4227 -37
rect -4139 -71 -4127 -37
rect -4239 -77 -4127 -71
rect -4061 -37 -3949 -31
rect -4061 -71 -4049 -37
rect -3961 -71 -3949 -37
rect -4061 -77 -3949 -71
rect -3883 -37 -3771 -31
rect -3883 -71 -3871 -37
rect -3783 -71 -3771 -37
rect -3883 -77 -3771 -71
rect -3705 -37 -3593 -31
rect -3705 -71 -3693 -37
rect -3605 -71 -3593 -37
rect -3705 -77 -3593 -71
rect -3527 -37 -3415 -31
rect -3527 -71 -3515 -37
rect -3427 -71 -3415 -37
rect -3527 -77 -3415 -71
rect -3349 -37 -3237 -31
rect -3349 -71 -3337 -37
rect -3249 -71 -3237 -37
rect -3349 -77 -3237 -71
rect -3171 -37 -3059 -31
rect -3171 -71 -3159 -37
rect -3071 -71 -3059 -37
rect -3171 -77 -3059 -71
rect -2993 -37 -2881 -31
rect -2993 -71 -2981 -37
rect -2893 -71 -2881 -37
rect -2993 -77 -2881 -71
rect -2815 -37 -2703 -31
rect -2815 -71 -2803 -37
rect -2715 -71 -2703 -37
rect -2815 -77 -2703 -71
rect -2637 -37 -2525 -31
rect -2637 -71 -2625 -37
rect -2537 -71 -2525 -37
rect -2637 -77 -2525 -71
rect -2459 -37 -2347 -31
rect -2459 -71 -2447 -37
rect -2359 -71 -2347 -37
rect -2459 -77 -2347 -71
rect -2281 -37 -2169 -31
rect -2281 -71 -2269 -37
rect -2181 -71 -2169 -37
rect -2281 -77 -2169 -71
rect -2103 -37 -1991 -31
rect -2103 -71 -2091 -37
rect -2003 -71 -1991 -37
rect -2103 -77 -1991 -71
rect -1925 -37 -1813 -31
rect -1925 -71 -1913 -37
rect -1825 -71 -1813 -37
rect -1925 -77 -1813 -71
rect -1747 -37 -1635 -31
rect -1747 -71 -1735 -37
rect -1647 -71 -1635 -37
rect -1747 -77 -1635 -71
rect -1569 -37 -1457 -31
rect -1569 -71 -1557 -37
rect -1469 -71 -1457 -37
rect -1569 -77 -1457 -71
rect -1391 -37 -1279 -31
rect -1391 -71 -1379 -37
rect -1291 -71 -1279 -37
rect -1391 -77 -1279 -71
rect -1213 -37 -1101 -31
rect -1213 -71 -1201 -37
rect -1113 -71 -1101 -37
rect -1213 -77 -1101 -71
rect -1035 -37 -923 -31
rect -1035 -71 -1023 -37
rect -935 -71 -923 -37
rect -1035 -77 -923 -71
rect -857 -37 -745 -31
rect -857 -71 -845 -37
rect -757 -71 -745 -37
rect -857 -77 -745 -71
rect -679 -37 -567 -31
rect -679 -71 -667 -37
rect -579 -71 -567 -37
rect -679 -77 -567 -71
rect -501 -37 -389 -31
rect -501 -71 -489 -37
rect -401 -71 -389 -37
rect -501 -77 -389 -71
rect -323 -37 -211 -31
rect -323 -71 -311 -37
rect -223 -71 -211 -37
rect -323 -77 -211 -71
rect -145 -37 -33 -31
rect -145 -71 -133 -37
rect -45 -71 -33 -37
rect -145 -77 -33 -71
rect 33 -37 145 -31
rect 33 -71 45 -37
rect 133 -71 145 -37
rect 33 -77 145 -71
rect 211 -37 323 -31
rect 211 -71 223 -37
rect 311 -71 323 -37
rect 211 -77 323 -71
rect 389 -37 501 -31
rect 389 -71 401 -37
rect 489 -71 501 -37
rect 389 -77 501 -71
rect 567 -37 679 -31
rect 567 -71 579 -37
rect 667 -71 679 -37
rect 567 -77 679 -71
rect 745 -37 857 -31
rect 745 -71 757 -37
rect 845 -71 857 -37
rect 745 -77 857 -71
rect 923 -37 1035 -31
rect 923 -71 935 -37
rect 1023 -71 1035 -37
rect 923 -77 1035 -71
rect 1101 -37 1213 -31
rect 1101 -71 1113 -37
rect 1201 -71 1213 -37
rect 1101 -77 1213 -71
rect 1279 -37 1391 -31
rect 1279 -71 1291 -37
rect 1379 -71 1391 -37
rect 1279 -77 1391 -71
rect 1457 -37 1569 -31
rect 1457 -71 1469 -37
rect 1557 -71 1569 -37
rect 1457 -77 1569 -71
rect 1635 -37 1747 -31
rect 1635 -71 1647 -37
rect 1735 -71 1747 -37
rect 1635 -77 1747 -71
rect 1813 -37 1925 -31
rect 1813 -71 1825 -37
rect 1913 -71 1925 -37
rect 1813 -77 1925 -71
rect 1991 -37 2103 -31
rect 1991 -71 2003 -37
rect 2091 -71 2103 -37
rect 1991 -77 2103 -71
rect 2169 -37 2281 -31
rect 2169 -71 2181 -37
rect 2269 -71 2281 -37
rect 2169 -77 2281 -71
rect 2347 -37 2459 -31
rect 2347 -71 2359 -37
rect 2447 -71 2459 -37
rect 2347 -77 2459 -71
rect 2525 -37 2637 -31
rect 2525 -71 2537 -37
rect 2625 -71 2637 -37
rect 2525 -77 2637 -71
rect 2703 -37 2815 -31
rect 2703 -71 2715 -37
rect 2803 -71 2815 -37
rect 2703 -77 2815 -71
rect 2881 -37 2993 -31
rect 2881 -71 2893 -37
rect 2981 -71 2993 -37
rect 2881 -77 2993 -71
rect 3059 -37 3171 -31
rect 3059 -71 3071 -37
rect 3159 -71 3171 -37
rect 3059 -77 3171 -71
rect 3237 -37 3349 -31
rect 3237 -71 3249 -37
rect 3337 -71 3349 -37
rect 3237 -77 3349 -71
rect 3415 -37 3527 -31
rect 3415 -71 3427 -37
rect 3515 -71 3527 -37
rect 3415 -77 3527 -71
rect 3593 -37 3705 -31
rect 3593 -71 3605 -37
rect 3693 -71 3705 -37
rect 3593 -77 3705 -71
rect 3771 -37 3883 -31
rect 3771 -71 3783 -37
rect 3871 -71 3883 -37
rect 3771 -77 3883 -71
rect 3949 -37 4061 -31
rect 3949 -71 3961 -37
rect 4049 -71 4061 -37
rect 3949 -77 4061 -71
rect 4127 -37 4239 -31
rect 4127 -71 4139 -37
rect 4227 -71 4239 -37
rect 4127 -77 4239 -71
rect 4305 -37 4417 -31
rect 4305 -71 4317 -37
rect 4405 -71 4417 -37
rect 4305 -77 4417 -71
rect 4483 -37 4595 -31
rect 4483 -71 4495 -37
rect 4583 -71 4595 -37
rect 4483 -77 4595 -71
rect 4661 -37 4773 -31
rect 4661 -71 4673 -37
rect 4761 -71 4773 -37
rect 4661 -77 4773 -71
rect 4839 -37 4951 -31
rect 4839 -71 4851 -37
rect 4939 -71 4951 -37
rect 4839 -77 4951 -71
rect 5017 -37 5129 -31
rect 5017 -71 5029 -37
rect 5117 -71 5129 -37
rect 5017 -77 5129 -71
rect 5195 -37 5307 -31
rect 5195 -71 5207 -37
rect 5295 -71 5307 -37
rect 5195 -77 5307 -71
rect 5373 -37 5485 -31
rect 5373 -71 5385 -37
rect 5473 -71 5485 -37
rect 5373 -77 5485 -71
rect 5551 -37 5663 -31
rect 5551 -71 5563 -37
rect 5651 -71 5663 -37
rect 5551 -77 5663 -71
rect 5729 -37 5841 -31
rect 5729 -71 5741 -37
rect 5829 -71 5841 -37
rect 5729 -77 5841 -71
rect 5907 -37 6019 -31
rect 5907 -71 5919 -37
rect 6007 -71 6019 -37
rect 5907 -77 6019 -71
rect 6085 -37 6197 -31
rect 6085 -71 6097 -37
rect 6185 -71 6197 -37
rect 6085 -77 6197 -71
rect 6263 -37 6375 -31
rect 6263 -71 6275 -37
rect 6363 -71 6375 -37
rect 6263 -77 6375 -71
rect 6441 -37 6553 -31
rect 6441 -71 6453 -37
rect 6541 -71 6553 -37
rect 6441 -77 6553 -71
rect 6619 -37 6731 -31
rect 6619 -71 6631 -37
rect 6719 -71 6731 -37
rect 6619 -77 6731 -71
rect 6797 -37 6909 -31
rect 6797 -71 6809 -37
rect 6897 -71 6909 -37
rect 6797 -77 6909 -71
rect 6975 -37 7087 -31
rect 6975 -71 6987 -37
rect 7075 -71 7087 -37
rect 6975 -77 7087 -71
rect 7153 -37 7265 -31
rect 7153 -71 7165 -37
rect 7253 -71 7265 -37
rect 7153 -77 7265 -71
rect 7331 -37 7443 -31
rect 7331 -71 7343 -37
rect 7431 -71 7443 -37
rect 7331 -77 7443 -71
rect 7509 -37 7621 -31
rect 7509 -71 7521 -37
rect 7609 -71 7621 -37
rect 7509 -77 7621 -71
rect 7687 -37 7799 -31
rect 7687 -71 7699 -37
rect 7787 -71 7799 -37
rect 7687 -77 7799 -71
rect 7865 -37 7977 -31
rect 7865 -71 7877 -37
rect 7965 -71 7977 -37
rect 7865 -77 7977 -71
rect -8033 -130 -7987 -118
rect -8033 -1306 -8027 -130
rect -7993 -1306 -7987 -130
rect -8033 -1318 -7987 -1306
rect -7855 -130 -7809 -118
rect -7855 -1306 -7849 -130
rect -7815 -1306 -7809 -130
rect -7855 -1318 -7809 -1306
rect -7677 -130 -7631 -118
rect -7677 -1306 -7671 -130
rect -7637 -1306 -7631 -130
rect -7677 -1318 -7631 -1306
rect -7499 -130 -7453 -118
rect -7499 -1306 -7493 -130
rect -7459 -1306 -7453 -130
rect -7499 -1318 -7453 -1306
rect -7321 -130 -7275 -118
rect -7321 -1306 -7315 -130
rect -7281 -1306 -7275 -130
rect -7321 -1318 -7275 -1306
rect -7143 -130 -7097 -118
rect -7143 -1306 -7137 -130
rect -7103 -1306 -7097 -130
rect -7143 -1318 -7097 -1306
rect -6965 -130 -6919 -118
rect -6965 -1306 -6959 -130
rect -6925 -1306 -6919 -130
rect -6965 -1318 -6919 -1306
rect -6787 -130 -6741 -118
rect -6787 -1306 -6781 -130
rect -6747 -1306 -6741 -130
rect -6787 -1318 -6741 -1306
rect -6609 -130 -6563 -118
rect -6609 -1306 -6603 -130
rect -6569 -1306 -6563 -130
rect -6609 -1318 -6563 -1306
rect -6431 -130 -6385 -118
rect -6431 -1306 -6425 -130
rect -6391 -1306 -6385 -130
rect -6431 -1318 -6385 -1306
rect -6253 -130 -6207 -118
rect -6253 -1306 -6247 -130
rect -6213 -1306 -6207 -130
rect -6253 -1318 -6207 -1306
rect -6075 -130 -6029 -118
rect -6075 -1306 -6069 -130
rect -6035 -1306 -6029 -130
rect -6075 -1318 -6029 -1306
rect -5897 -130 -5851 -118
rect -5897 -1306 -5891 -130
rect -5857 -1306 -5851 -130
rect -5897 -1318 -5851 -1306
rect -5719 -130 -5673 -118
rect -5719 -1306 -5713 -130
rect -5679 -1306 -5673 -130
rect -5719 -1318 -5673 -1306
rect -5541 -130 -5495 -118
rect -5541 -1306 -5535 -130
rect -5501 -1306 -5495 -130
rect -5541 -1318 -5495 -1306
rect -5363 -130 -5317 -118
rect -5363 -1306 -5357 -130
rect -5323 -1306 -5317 -130
rect -5363 -1318 -5317 -1306
rect -5185 -130 -5139 -118
rect -5185 -1306 -5179 -130
rect -5145 -1306 -5139 -130
rect -5185 -1318 -5139 -1306
rect -5007 -130 -4961 -118
rect -5007 -1306 -5001 -130
rect -4967 -1306 -4961 -130
rect -5007 -1318 -4961 -1306
rect -4829 -130 -4783 -118
rect -4829 -1306 -4823 -130
rect -4789 -1306 -4783 -130
rect -4829 -1318 -4783 -1306
rect -4651 -130 -4605 -118
rect -4651 -1306 -4645 -130
rect -4611 -1306 -4605 -130
rect -4651 -1318 -4605 -1306
rect -4473 -130 -4427 -118
rect -4473 -1306 -4467 -130
rect -4433 -1306 -4427 -130
rect -4473 -1318 -4427 -1306
rect -4295 -130 -4249 -118
rect -4295 -1306 -4289 -130
rect -4255 -1306 -4249 -130
rect -4295 -1318 -4249 -1306
rect -4117 -130 -4071 -118
rect -4117 -1306 -4111 -130
rect -4077 -1306 -4071 -130
rect -4117 -1318 -4071 -1306
rect -3939 -130 -3893 -118
rect -3939 -1306 -3933 -130
rect -3899 -1306 -3893 -130
rect -3939 -1318 -3893 -1306
rect -3761 -130 -3715 -118
rect -3761 -1306 -3755 -130
rect -3721 -1306 -3715 -130
rect -3761 -1318 -3715 -1306
rect -3583 -130 -3537 -118
rect -3583 -1306 -3577 -130
rect -3543 -1306 -3537 -130
rect -3583 -1318 -3537 -1306
rect -3405 -130 -3359 -118
rect -3405 -1306 -3399 -130
rect -3365 -1306 -3359 -130
rect -3405 -1318 -3359 -1306
rect -3227 -130 -3181 -118
rect -3227 -1306 -3221 -130
rect -3187 -1306 -3181 -130
rect -3227 -1318 -3181 -1306
rect -3049 -130 -3003 -118
rect -3049 -1306 -3043 -130
rect -3009 -1306 -3003 -130
rect -3049 -1318 -3003 -1306
rect -2871 -130 -2825 -118
rect -2871 -1306 -2865 -130
rect -2831 -1306 -2825 -130
rect -2871 -1318 -2825 -1306
rect -2693 -130 -2647 -118
rect -2693 -1306 -2687 -130
rect -2653 -1306 -2647 -130
rect -2693 -1318 -2647 -1306
rect -2515 -130 -2469 -118
rect -2515 -1306 -2509 -130
rect -2475 -1306 -2469 -130
rect -2515 -1318 -2469 -1306
rect -2337 -130 -2291 -118
rect -2337 -1306 -2331 -130
rect -2297 -1306 -2291 -130
rect -2337 -1318 -2291 -1306
rect -2159 -130 -2113 -118
rect -2159 -1306 -2153 -130
rect -2119 -1306 -2113 -130
rect -2159 -1318 -2113 -1306
rect -1981 -130 -1935 -118
rect -1981 -1306 -1975 -130
rect -1941 -1306 -1935 -130
rect -1981 -1318 -1935 -1306
rect -1803 -130 -1757 -118
rect -1803 -1306 -1797 -130
rect -1763 -1306 -1757 -130
rect -1803 -1318 -1757 -1306
rect -1625 -130 -1579 -118
rect -1625 -1306 -1619 -130
rect -1585 -1306 -1579 -130
rect -1625 -1318 -1579 -1306
rect -1447 -130 -1401 -118
rect -1447 -1306 -1441 -130
rect -1407 -1306 -1401 -130
rect -1447 -1318 -1401 -1306
rect -1269 -130 -1223 -118
rect -1269 -1306 -1263 -130
rect -1229 -1306 -1223 -130
rect -1269 -1318 -1223 -1306
rect -1091 -130 -1045 -118
rect -1091 -1306 -1085 -130
rect -1051 -1306 -1045 -130
rect -1091 -1318 -1045 -1306
rect -913 -130 -867 -118
rect -913 -1306 -907 -130
rect -873 -1306 -867 -130
rect -913 -1318 -867 -1306
rect -735 -130 -689 -118
rect -735 -1306 -729 -130
rect -695 -1306 -689 -130
rect -735 -1318 -689 -1306
rect -557 -130 -511 -118
rect -557 -1306 -551 -130
rect -517 -1306 -511 -130
rect -557 -1318 -511 -1306
rect -379 -130 -333 -118
rect -379 -1306 -373 -130
rect -339 -1306 -333 -130
rect -379 -1318 -333 -1306
rect -201 -130 -155 -118
rect -201 -1306 -195 -130
rect -161 -1306 -155 -130
rect -201 -1318 -155 -1306
rect -23 -130 23 -118
rect -23 -1306 -17 -130
rect 17 -1306 23 -130
rect -23 -1318 23 -1306
rect 155 -130 201 -118
rect 155 -1306 161 -130
rect 195 -1306 201 -130
rect 155 -1318 201 -1306
rect 333 -130 379 -118
rect 333 -1306 339 -130
rect 373 -1306 379 -130
rect 333 -1318 379 -1306
rect 511 -130 557 -118
rect 511 -1306 517 -130
rect 551 -1306 557 -130
rect 511 -1318 557 -1306
rect 689 -130 735 -118
rect 689 -1306 695 -130
rect 729 -1306 735 -130
rect 689 -1318 735 -1306
rect 867 -130 913 -118
rect 867 -1306 873 -130
rect 907 -1306 913 -130
rect 867 -1318 913 -1306
rect 1045 -130 1091 -118
rect 1045 -1306 1051 -130
rect 1085 -1306 1091 -130
rect 1045 -1318 1091 -1306
rect 1223 -130 1269 -118
rect 1223 -1306 1229 -130
rect 1263 -1306 1269 -130
rect 1223 -1318 1269 -1306
rect 1401 -130 1447 -118
rect 1401 -1306 1407 -130
rect 1441 -1306 1447 -130
rect 1401 -1318 1447 -1306
rect 1579 -130 1625 -118
rect 1579 -1306 1585 -130
rect 1619 -1306 1625 -130
rect 1579 -1318 1625 -1306
rect 1757 -130 1803 -118
rect 1757 -1306 1763 -130
rect 1797 -1306 1803 -130
rect 1757 -1318 1803 -1306
rect 1935 -130 1981 -118
rect 1935 -1306 1941 -130
rect 1975 -1306 1981 -130
rect 1935 -1318 1981 -1306
rect 2113 -130 2159 -118
rect 2113 -1306 2119 -130
rect 2153 -1306 2159 -130
rect 2113 -1318 2159 -1306
rect 2291 -130 2337 -118
rect 2291 -1306 2297 -130
rect 2331 -1306 2337 -130
rect 2291 -1318 2337 -1306
rect 2469 -130 2515 -118
rect 2469 -1306 2475 -130
rect 2509 -1306 2515 -130
rect 2469 -1318 2515 -1306
rect 2647 -130 2693 -118
rect 2647 -1306 2653 -130
rect 2687 -1306 2693 -130
rect 2647 -1318 2693 -1306
rect 2825 -130 2871 -118
rect 2825 -1306 2831 -130
rect 2865 -1306 2871 -130
rect 2825 -1318 2871 -1306
rect 3003 -130 3049 -118
rect 3003 -1306 3009 -130
rect 3043 -1306 3049 -130
rect 3003 -1318 3049 -1306
rect 3181 -130 3227 -118
rect 3181 -1306 3187 -130
rect 3221 -1306 3227 -130
rect 3181 -1318 3227 -1306
rect 3359 -130 3405 -118
rect 3359 -1306 3365 -130
rect 3399 -1306 3405 -130
rect 3359 -1318 3405 -1306
rect 3537 -130 3583 -118
rect 3537 -1306 3543 -130
rect 3577 -1306 3583 -130
rect 3537 -1318 3583 -1306
rect 3715 -130 3761 -118
rect 3715 -1306 3721 -130
rect 3755 -1306 3761 -130
rect 3715 -1318 3761 -1306
rect 3893 -130 3939 -118
rect 3893 -1306 3899 -130
rect 3933 -1306 3939 -130
rect 3893 -1318 3939 -1306
rect 4071 -130 4117 -118
rect 4071 -1306 4077 -130
rect 4111 -1306 4117 -130
rect 4071 -1318 4117 -1306
rect 4249 -130 4295 -118
rect 4249 -1306 4255 -130
rect 4289 -1306 4295 -130
rect 4249 -1318 4295 -1306
rect 4427 -130 4473 -118
rect 4427 -1306 4433 -130
rect 4467 -1306 4473 -130
rect 4427 -1318 4473 -1306
rect 4605 -130 4651 -118
rect 4605 -1306 4611 -130
rect 4645 -1306 4651 -130
rect 4605 -1318 4651 -1306
rect 4783 -130 4829 -118
rect 4783 -1306 4789 -130
rect 4823 -1306 4829 -130
rect 4783 -1318 4829 -1306
rect 4961 -130 5007 -118
rect 4961 -1306 4967 -130
rect 5001 -1306 5007 -130
rect 4961 -1318 5007 -1306
rect 5139 -130 5185 -118
rect 5139 -1306 5145 -130
rect 5179 -1306 5185 -130
rect 5139 -1318 5185 -1306
rect 5317 -130 5363 -118
rect 5317 -1306 5323 -130
rect 5357 -1306 5363 -130
rect 5317 -1318 5363 -1306
rect 5495 -130 5541 -118
rect 5495 -1306 5501 -130
rect 5535 -1306 5541 -130
rect 5495 -1318 5541 -1306
rect 5673 -130 5719 -118
rect 5673 -1306 5679 -130
rect 5713 -1306 5719 -130
rect 5673 -1318 5719 -1306
rect 5851 -130 5897 -118
rect 5851 -1306 5857 -130
rect 5891 -1306 5897 -130
rect 5851 -1318 5897 -1306
rect 6029 -130 6075 -118
rect 6029 -1306 6035 -130
rect 6069 -1306 6075 -130
rect 6029 -1318 6075 -1306
rect 6207 -130 6253 -118
rect 6207 -1306 6213 -130
rect 6247 -1306 6253 -130
rect 6207 -1318 6253 -1306
rect 6385 -130 6431 -118
rect 6385 -1306 6391 -130
rect 6425 -1306 6431 -130
rect 6385 -1318 6431 -1306
rect 6563 -130 6609 -118
rect 6563 -1306 6569 -130
rect 6603 -1306 6609 -130
rect 6563 -1318 6609 -1306
rect 6741 -130 6787 -118
rect 6741 -1306 6747 -130
rect 6781 -1306 6787 -130
rect 6741 -1318 6787 -1306
rect 6919 -130 6965 -118
rect 6919 -1306 6925 -130
rect 6959 -1306 6965 -130
rect 6919 -1318 6965 -1306
rect 7097 -130 7143 -118
rect 7097 -1306 7103 -130
rect 7137 -1306 7143 -130
rect 7097 -1318 7143 -1306
rect 7275 -130 7321 -118
rect 7275 -1306 7281 -130
rect 7315 -1306 7321 -130
rect 7275 -1318 7321 -1306
rect 7453 -130 7499 -118
rect 7453 -1306 7459 -130
rect 7493 -1306 7499 -130
rect 7453 -1318 7499 -1306
rect 7631 -130 7677 -118
rect 7631 -1306 7637 -130
rect 7671 -1306 7677 -130
rect 7631 -1318 7677 -1306
rect 7809 -130 7855 -118
rect 7809 -1306 7815 -130
rect 7849 -1306 7855 -130
rect 7809 -1318 7855 -1306
rect 7987 -130 8033 -118
rect 7987 -1306 7993 -130
rect 8027 -1306 8033 -130
rect 7987 -1318 8033 -1306
rect -7977 -1365 -7865 -1359
rect -7977 -1399 -7965 -1365
rect -7877 -1399 -7865 -1365
rect -7977 -1405 -7865 -1399
rect -7799 -1365 -7687 -1359
rect -7799 -1399 -7787 -1365
rect -7699 -1399 -7687 -1365
rect -7799 -1405 -7687 -1399
rect -7621 -1365 -7509 -1359
rect -7621 -1399 -7609 -1365
rect -7521 -1399 -7509 -1365
rect -7621 -1405 -7509 -1399
rect -7443 -1365 -7331 -1359
rect -7443 -1399 -7431 -1365
rect -7343 -1399 -7331 -1365
rect -7443 -1405 -7331 -1399
rect -7265 -1365 -7153 -1359
rect -7265 -1399 -7253 -1365
rect -7165 -1399 -7153 -1365
rect -7265 -1405 -7153 -1399
rect -7087 -1365 -6975 -1359
rect -7087 -1399 -7075 -1365
rect -6987 -1399 -6975 -1365
rect -7087 -1405 -6975 -1399
rect -6909 -1365 -6797 -1359
rect -6909 -1399 -6897 -1365
rect -6809 -1399 -6797 -1365
rect -6909 -1405 -6797 -1399
rect -6731 -1365 -6619 -1359
rect -6731 -1399 -6719 -1365
rect -6631 -1399 -6619 -1365
rect -6731 -1405 -6619 -1399
rect -6553 -1365 -6441 -1359
rect -6553 -1399 -6541 -1365
rect -6453 -1399 -6441 -1365
rect -6553 -1405 -6441 -1399
rect -6375 -1365 -6263 -1359
rect -6375 -1399 -6363 -1365
rect -6275 -1399 -6263 -1365
rect -6375 -1405 -6263 -1399
rect -6197 -1365 -6085 -1359
rect -6197 -1399 -6185 -1365
rect -6097 -1399 -6085 -1365
rect -6197 -1405 -6085 -1399
rect -6019 -1365 -5907 -1359
rect -6019 -1399 -6007 -1365
rect -5919 -1399 -5907 -1365
rect -6019 -1405 -5907 -1399
rect -5841 -1365 -5729 -1359
rect -5841 -1399 -5829 -1365
rect -5741 -1399 -5729 -1365
rect -5841 -1405 -5729 -1399
rect -5663 -1365 -5551 -1359
rect -5663 -1399 -5651 -1365
rect -5563 -1399 -5551 -1365
rect -5663 -1405 -5551 -1399
rect -5485 -1365 -5373 -1359
rect -5485 -1399 -5473 -1365
rect -5385 -1399 -5373 -1365
rect -5485 -1405 -5373 -1399
rect -5307 -1365 -5195 -1359
rect -5307 -1399 -5295 -1365
rect -5207 -1399 -5195 -1365
rect -5307 -1405 -5195 -1399
rect -5129 -1365 -5017 -1359
rect -5129 -1399 -5117 -1365
rect -5029 -1399 -5017 -1365
rect -5129 -1405 -5017 -1399
rect -4951 -1365 -4839 -1359
rect -4951 -1399 -4939 -1365
rect -4851 -1399 -4839 -1365
rect -4951 -1405 -4839 -1399
rect -4773 -1365 -4661 -1359
rect -4773 -1399 -4761 -1365
rect -4673 -1399 -4661 -1365
rect -4773 -1405 -4661 -1399
rect -4595 -1365 -4483 -1359
rect -4595 -1399 -4583 -1365
rect -4495 -1399 -4483 -1365
rect -4595 -1405 -4483 -1399
rect -4417 -1365 -4305 -1359
rect -4417 -1399 -4405 -1365
rect -4317 -1399 -4305 -1365
rect -4417 -1405 -4305 -1399
rect -4239 -1365 -4127 -1359
rect -4239 -1399 -4227 -1365
rect -4139 -1399 -4127 -1365
rect -4239 -1405 -4127 -1399
rect -4061 -1365 -3949 -1359
rect -4061 -1399 -4049 -1365
rect -3961 -1399 -3949 -1365
rect -4061 -1405 -3949 -1399
rect -3883 -1365 -3771 -1359
rect -3883 -1399 -3871 -1365
rect -3783 -1399 -3771 -1365
rect -3883 -1405 -3771 -1399
rect -3705 -1365 -3593 -1359
rect -3705 -1399 -3693 -1365
rect -3605 -1399 -3593 -1365
rect -3705 -1405 -3593 -1399
rect -3527 -1365 -3415 -1359
rect -3527 -1399 -3515 -1365
rect -3427 -1399 -3415 -1365
rect -3527 -1405 -3415 -1399
rect -3349 -1365 -3237 -1359
rect -3349 -1399 -3337 -1365
rect -3249 -1399 -3237 -1365
rect -3349 -1405 -3237 -1399
rect -3171 -1365 -3059 -1359
rect -3171 -1399 -3159 -1365
rect -3071 -1399 -3059 -1365
rect -3171 -1405 -3059 -1399
rect -2993 -1365 -2881 -1359
rect -2993 -1399 -2981 -1365
rect -2893 -1399 -2881 -1365
rect -2993 -1405 -2881 -1399
rect -2815 -1365 -2703 -1359
rect -2815 -1399 -2803 -1365
rect -2715 -1399 -2703 -1365
rect -2815 -1405 -2703 -1399
rect -2637 -1365 -2525 -1359
rect -2637 -1399 -2625 -1365
rect -2537 -1399 -2525 -1365
rect -2637 -1405 -2525 -1399
rect -2459 -1365 -2347 -1359
rect -2459 -1399 -2447 -1365
rect -2359 -1399 -2347 -1365
rect -2459 -1405 -2347 -1399
rect -2281 -1365 -2169 -1359
rect -2281 -1399 -2269 -1365
rect -2181 -1399 -2169 -1365
rect -2281 -1405 -2169 -1399
rect -2103 -1365 -1991 -1359
rect -2103 -1399 -2091 -1365
rect -2003 -1399 -1991 -1365
rect -2103 -1405 -1991 -1399
rect -1925 -1365 -1813 -1359
rect -1925 -1399 -1913 -1365
rect -1825 -1399 -1813 -1365
rect -1925 -1405 -1813 -1399
rect -1747 -1365 -1635 -1359
rect -1747 -1399 -1735 -1365
rect -1647 -1399 -1635 -1365
rect -1747 -1405 -1635 -1399
rect -1569 -1365 -1457 -1359
rect -1569 -1399 -1557 -1365
rect -1469 -1399 -1457 -1365
rect -1569 -1405 -1457 -1399
rect -1391 -1365 -1279 -1359
rect -1391 -1399 -1379 -1365
rect -1291 -1399 -1279 -1365
rect -1391 -1405 -1279 -1399
rect -1213 -1365 -1101 -1359
rect -1213 -1399 -1201 -1365
rect -1113 -1399 -1101 -1365
rect -1213 -1405 -1101 -1399
rect -1035 -1365 -923 -1359
rect -1035 -1399 -1023 -1365
rect -935 -1399 -923 -1365
rect -1035 -1405 -923 -1399
rect -857 -1365 -745 -1359
rect -857 -1399 -845 -1365
rect -757 -1399 -745 -1365
rect -857 -1405 -745 -1399
rect -679 -1365 -567 -1359
rect -679 -1399 -667 -1365
rect -579 -1399 -567 -1365
rect -679 -1405 -567 -1399
rect -501 -1365 -389 -1359
rect -501 -1399 -489 -1365
rect -401 -1399 -389 -1365
rect -501 -1405 -389 -1399
rect -323 -1365 -211 -1359
rect -323 -1399 -311 -1365
rect -223 -1399 -211 -1365
rect -323 -1405 -211 -1399
rect -145 -1365 -33 -1359
rect -145 -1399 -133 -1365
rect -45 -1399 -33 -1365
rect -145 -1405 -33 -1399
rect 33 -1365 145 -1359
rect 33 -1399 45 -1365
rect 133 -1399 145 -1365
rect 33 -1405 145 -1399
rect 211 -1365 323 -1359
rect 211 -1399 223 -1365
rect 311 -1399 323 -1365
rect 211 -1405 323 -1399
rect 389 -1365 501 -1359
rect 389 -1399 401 -1365
rect 489 -1399 501 -1365
rect 389 -1405 501 -1399
rect 567 -1365 679 -1359
rect 567 -1399 579 -1365
rect 667 -1399 679 -1365
rect 567 -1405 679 -1399
rect 745 -1365 857 -1359
rect 745 -1399 757 -1365
rect 845 -1399 857 -1365
rect 745 -1405 857 -1399
rect 923 -1365 1035 -1359
rect 923 -1399 935 -1365
rect 1023 -1399 1035 -1365
rect 923 -1405 1035 -1399
rect 1101 -1365 1213 -1359
rect 1101 -1399 1113 -1365
rect 1201 -1399 1213 -1365
rect 1101 -1405 1213 -1399
rect 1279 -1365 1391 -1359
rect 1279 -1399 1291 -1365
rect 1379 -1399 1391 -1365
rect 1279 -1405 1391 -1399
rect 1457 -1365 1569 -1359
rect 1457 -1399 1469 -1365
rect 1557 -1399 1569 -1365
rect 1457 -1405 1569 -1399
rect 1635 -1365 1747 -1359
rect 1635 -1399 1647 -1365
rect 1735 -1399 1747 -1365
rect 1635 -1405 1747 -1399
rect 1813 -1365 1925 -1359
rect 1813 -1399 1825 -1365
rect 1913 -1399 1925 -1365
rect 1813 -1405 1925 -1399
rect 1991 -1365 2103 -1359
rect 1991 -1399 2003 -1365
rect 2091 -1399 2103 -1365
rect 1991 -1405 2103 -1399
rect 2169 -1365 2281 -1359
rect 2169 -1399 2181 -1365
rect 2269 -1399 2281 -1365
rect 2169 -1405 2281 -1399
rect 2347 -1365 2459 -1359
rect 2347 -1399 2359 -1365
rect 2447 -1399 2459 -1365
rect 2347 -1405 2459 -1399
rect 2525 -1365 2637 -1359
rect 2525 -1399 2537 -1365
rect 2625 -1399 2637 -1365
rect 2525 -1405 2637 -1399
rect 2703 -1365 2815 -1359
rect 2703 -1399 2715 -1365
rect 2803 -1399 2815 -1365
rect 2703 -1405 2815 -1399
rect 2881 -1365 2993 -1359
rect 2881 -1399 2893 -1365
rect 2981 -1399 2993 -1365
rect 2881 -1405 2993 -1399
rect 3059 -1365 3171 -1359
rect 3059 -1399 3071 -1365
rect 3159 -1399 3171 -1365
rect 3059 -1405 3171 -1399
rect 3237 -1365 3349 -1359
rect 3237 -1399 3249 -1365
rect 3337 -1399 3349 -1365
rect 3237 -1405 3349 -1399
rect 3415 -1365 3527 -1359
rect 3415 -1399 3427 -1365
rect 3515 -1399 3527 -1365
rect 3415 -1405 3527 -1399
rect 3593 -1365 3705 -1359
rect 3593 -1399 3605 -1365
rect 3693 -1399 3705 -1365
rect 3593 -1405 3705 -1399
rect 3771 -1365 3883 -1359
rect 3771 -1399 3783 -1365
rect 3871 -1399 3883 -1365
rect 3771 -1405 3883 -1399
rect 3949 -1365 4061 -1359
rect 3949 -1399 3961 -1365
rect 4049 -1399 4061 -1365
rect 3949 -1405 4061 -1399
rect 4127 -1365 4239 -1359
rect 4127 -1399 4139 -1365
rect 4227 -1399 4239 -1365
rect 4127 -1405 4239 -1399
rect 4305 -1365 4417 -1359
rect 4305 -1399 4317 -1365
rect 4405 -1399 4417 -1365
rect 4305 -1405 4417 -1399
rect 4483 -1365 4595 -1359
rect 4483 -1399 4495 -1365
rect 4583 -1399 4595 -1365
rect 4483 -1405 4595 -1399
rect 4661 -1365 4773 -1359
rect 4661 -1399 4673 -1365
rect 4761 -1399 4773 -1365
rect 4661 -1405 4773 -1399
rect 4839 -1365 4951 -1359
rect 4839 -1399 4851 -1365
rect 4939 -1399 4951 -1365
rect 4839 -1405 4951 -1399
rect 5017 -1365 5129 -1359
rect 5017 -1399 5029 -1365
rect 5117 -1399 5129 -1365
rect 5017 -1405 5129 -1399
rect 5195 -1365 5307 -1359
rect 5195 -1399 5207 -1365
rect 5295 -1399 5307 -1365
rect 5195 -1405 5307 -1399
rect 5373 -1365 5485 -1359
rect 5373 -1399 5385 -1365
rect 5473 -1399 5485 -1365
rect 5373 -1405 5485 -1399
rect 5551 -1365 5663 -1359
rect 5551 -1399 5563 -1365
rect 5651 -1399 5663 -1365
rect 5551 -1405 5663 -1399
rect 5729 -1365 5841 -1359
rect 5729 -1399 5741 -1365
rect 5829 -1399 5841 -1365
rect 5729 -1405 5841 -1399
rect 5907 -1365 6019 -1359
rect 5907 -1399 5919 -1365
rect 6007 -1399 6019 -1365
rect 5907 -1405 6019 -1399
rect 6085 -1365 6197 -1359
rect 6085 -1399 6097 -1365
rect 6185 -1399 6197 -1365
rect 6085 -1405 6197 -1399
rect 6263 -1365 6375 -1359
rect 6263 -1399 6275 -1365
rect 6363 -1399 6375 -1365
rect 6263 -1405 6375 -1399
rect 6441 -1365 6553 -1359
rect 6441 -1399 6453 -1365
rect 6541 -1399 6553 -1365
rect 6441 -1405 6553 -1399
rect 6619 -1365 6731 -1359
rect 6619 -1399 6631 -1365
rect 6719 -1399 6731 -1365
rect 6619 -1405 6731 -1399
rect 6797 -1365 6909 -1359
rect 6797 -1399 6809 -1365
rect 6897 -1399 6909 -1365
rect 6797 -1405 6909 -1399
rect 6975 -1365 7087 -1359
rect 6975 -1399 6987 -1365
rect 7075 -1399 7087 -1365
rect 6975 -1405 7087 -1399
rect 7153 -1365 7265 -1359
rect 7153 -1399 7165 -1365
rect 7253 -1399 7265 -1365
rect 7153 -1405 7265 -1399
rect 7331 -1365 7443 -1359
rect 7331 -1399 7343 -1365
rect 7431 -1399 7443 -1365
rect 7331 -1405 7443 -1399
rect 7509 -1365 7621 -1359
rect 7509 -1399 7521 -1365
rect 7609 -1399 7621 -1365
rect 7509 -1405 7621 -1399
rect 7687 -1365 7799 -1359
rect 7687 -1399 7699 -1365
rect 7787 -1399 7799 -1365
rect 7687 -1405 7799 -1399
rect 7865 -1365 7977 -1359
rect 7865 -1399 7877 -1365
rect 7965 -1399 7977 -1365
rect 7865 -1405 7977 -1399
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -8124 -1484 8124 1484
string parameters w 6 l 0.6 m 2 nf 90 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
