magic
tech sky130B
magscale 1 2
timestamp 1606423539
<< error_p >>
rect -2920 1635 -2862 1641
rect -2802 1635 -2744 1641
rect -2684 1635 -2626 1641
rect -2566 1635 -2508 1641
rect -2448 1635 -2390 1641
rect -2330 1635 -2272 1641
rect -2212 1635 -2154 1641
rect -2094 1635 -2036 1641
rect -1976 1635 -1918 1641
rect -1858 1635 -1800 1641
rect -1740 1635 -1682 1641
rect -1622 1635 -1564 1641
rect -1504 1635 -1446 1641
rect -1386 1635 -1328 1641
rect -1268 1635 -1210 1641
rect -1150 1635 -1092 1641
rect -1032 1635 -974 1641
rect -914 1635 -856 1641
rect -796 1635 -738 1641
rect -678 1635 -620 1641
rect -560 1635 -502 1641
rect -442 1635 -384 1641
rect -324 1635 -266 1641
rect -206 1635 -148 1641
rect -88 1635 -30 1641
rect 30 1635 88 1641
rect 148 1635 206 1641
rect 266 1635 324 1641
rect 384 1635 442 1641
rect 502 1635 560 1641
rect 620 1635 678 1641
rect 738 1635 796 1641
rect 856 1635 914 1641
rect 974 1635 1032 1641
rect 1092 1635 1150 1641
rect 1210 1635 1268 1641
rect 1328 1635 1386 1641
rect 1446 1635 1504 1641
rect 1564 1635 1622 1641
rect 1682 1635 1740 1641
rect 1800 1635 1858 1641
rect 1918 1635 1976 1641
rect 2036 1635 2094 1641
rect 2154 1635 2212 1641
rect 2272 1635 2330 1641
rect 2390 1635 2448 1641
rect 2508 1635 2566 1641
rect 2626 1635 2684 1641
rect 2744 1635 2802 1641
rect 2862 1635 2920 1641
rect -2920 1601 -2908 1635
rect -2802 1601 -2790 1635
rect -2684 1601 -2672 1635
rect -2566 1601 -2554 1635
rect -2448 1601 -2436 1635
rect -2330 1601 -2318 1635
rect -2212 1601 -2200 1635
rect -2094 1601 -2082 1635
rect -1976 1601 -1964 1635
rect -1858 1601 -1846 1635
rect -1740 1601 -1728 1635
rect -1622 1601 -1610 1635
rect -1504 1601 -1492 1635
rect -1386 1601 -1374 1635
rect -1268 1601 -1256 1635
rect -1150 1601 -1138 1635
rect -1032 1601 -1020 1635
rect -914 1601 -902 1635
rect -796 1601 -784 1635
rect -678 1601 -666 1635
rect -560 1601 -548 1635
rect -442 1601 -430 1635
rect -324 1601 -312 1635
rect -206 1601 -194 1635
rect -88 1601 -76 1635
rect 30 1601 42 1635
rect 148 1601 160 1635
rect 266 1601 278 1635
rect 384 1601 396 1635
rect 502 1601 514 1635
rect 620 1601 632 1635
rect 738 1601 750 1635
rect 856 1601 868 1635
rect 974 1601 986 1635
rect 1092 1601 1104 1635
rect 1210 1601 1222 1635
rect 1328 1601 1340 1635
rect 1446 1601 1458 1635
rect 1564 1601 1576 1635
rect 1682 1601 1694 1635
rect 1800 1601 1812 1635
rect 1918 1601 1930 1635
rect 2036 1601 2048 1635
rect 2154 1601 2166 1635
rect 2272 1601 2284 1635
rect 2390 1601 2402 1635
rect 2508 1601 2520 1635
rect 2626 1601 2638 1635
rect 2744 1601 2756 1635
rect 2862 1601 2874 1635
rect -2920 1595 -2862 1601
rect -2802 1595 -2744 1601
rect -2684 1595 -2626 1601
rect -2566 1595 -2508 1601
rect -2448 1595 -2390 1601
rect -2330 1595 -2272 1601
rect -2212 1595 -2154 1601
rect -2094 1595 -2036 1601
rect -1976 1595 -1918 1601
rect -1858 1595 -1800 1601
rect -1740 1595 -1682 1601
rect -1622 1595 -1564 1601
rect -1504 1595 -1446 1601
rect -1386 1595 -1328 1601
rect -1268 1595 -1210 1601
rect -1150 1595 -1092 1601
rect -1032 1595 -974 1601
rect -914 1595 -856 1601
rect -796 1595 -738 1601
rect -678 1595 -620 1601
rect -560 1595 -502 1601
rect -442 1595 -384 1601
rect -324 1595 -266 1601
rect -206 1595 -148 1601
rect -88 1595 -30 1601
rect 30 1595 88 1601
rect 148 1595 206 1601
rect 266 1595 324 1601
rect 384 1595 442 1601
rect 502 1595 560 1601
rect 620 1595 678 1601
rect 738 1595 796 1601
rect 856 1595 914 1601
rect 974 1595 1032 1601
rect 1092 1595 1150 1601
rect 1210 1595 1268 1601
rect 1328 1595 1386 1601
rect 1446 1595 1504 1601
rect 1564 1595 1622 1601
rect 1682 1595 1740 1601
rect 1800 1595 1858 1601
rect 1918 1595 1976 1601
rect 2036 1595 2094 1601
rect 2154 1595 2212 1601
rect 2272 1595 2330 1601
rect 2390 1595 2448 1601
rect 2508 1595 2566 1601
rect 2626 1595 2684 1601
rect 2744 1595 2802 1601
rect 2862 1595 2920 1601
rect -2920 907 -2862 913
rect -2802 907 -2744 913
rect -2684 907 -2626 913
rect -2566 907 -2508 913
rect -2448 907 -2390 913
rect -2330 907 -2272 913
rect -2212 907 -2154 913
rect -2094 907 -2036 913
rect -1976 907 -1918 913
rect -1858 907 -1800 913
rect -1740 907 -1682 913
rect -1622 907 -1564 913
rect -1504 907 -1446 913
rect -1386 907 -1328 913
rect -1268 907 -1210 913
rect -1150 907 -1092 913
rect -1032 907 -974 913
rect -914 907 -856 913
rect -796 907 -738 913
rect -678 907 -620 913
rect -560 907 -502 913
rect -442 907 -384 913
rect -324 907 -266 913
rect -206 907 -148 913
rect -88 907 -30 913
rect 30 907 88 913
rect 148 907 206 913
rect 266 907 324 913
rect 384 907 442 913
rect 502 907 560 913
rect 620 907 678 913
rect 738 907 796 913
rect 856 907 914 913
rect 974 907 1032 913
rect 1092 907 1150 913
rect 1210 907 1268 913
rect 1328 907 1386 913
rect 1446 907 1504 913
rect 1564 907 1622 913
rect 1682 907 1740 913
rect 1800 907 1858 913
rect 1918 907 1976 913
rect 2036 907 2094 913
rect 2154 907 2212 913
rect 2272 907 2330 913
rect 2390 907 2448 913
rect 2508 907 2566 913
rect 2626 907 2684 913
rect 2744 907 2802 913
rect 2862 907 2920 913
rect -2920 873 -2908 907
rect -2802 873 -2790 907
rect -2684 873 -2672 907
rect -2566 873 -2554 907
rect -2448 873 -2436 907
rect -2330 873 -2318 907
rect -2212 873 -2200 907
rect -2094 873 -2082 907
rect -1976 873 -1964 907
rect -1858 873 -1846 907
rect -1740 873 -1728 907
rect -1622 873 -1610 907
rect -1504 873 -1492 907
rect -1386 873 -1374 907
rect -1268 873 -1256 907
rect -1150 873 -1138 907
rect -1032 873 -1020 907
rect -914 873 -902 907
rect -796 873 -784 907
rect -678 873 -666 907
rect -560 873 -548 907
rect -442 873 -430 907
rect -324 873 -312 907
rect -206 873 -194 907
rect -88 873 -76 907
rect 30 873 42 907
rect 148 873 160 907
rect 266 873 278 907
rect 384 873 396 907
rect 502 873 514 907
rect 620 873 632 907
rect 738 873 750 907
rect 856 873 868 907
rect 974 873 986 907
rect 1092 873 1104 907
rect 1210 873 1222 907
rect 1328 873 1340 907
rect 1446 873 1458 907
rect 1564 873 1576 907
rect 1682 873 1694 907
rect 1800 873 1812 907
rect 1918 873 1930 907
rect 2036 873 2048 907
rect 2154 873 2166 907
rect 2272 873 2284 907
rect 2390 873 2402 907
rect 2508 873 2520 907
rect 2626 873 2638 907
rect 2744 873 2756 907
rect 2862 873 2874 907
rect -2920 867 -2862 873
rect -2802 867 -2744 873
rect -2684 867 -2626 873
rect -2566 867 -2508 873
rect -2448 867 -2390 873
rect -2330 867 -2272 873
rect -2212 867 -2154 873
rect -2094 867 -2036 873
rect -1976 867 -1918 873
rect -1858 867 -1800 873
rect -1740 867 -1682 873
rect -1622 867 -1564 873
rect -1504 867 -1446 873
rect -1386 867 -1328 873
rect -1268 867 -1210 873
rect -1150 867 -1092 873
rect -1032 867 -974 873
rect -914 867 -856 873
rect -796 867 -738 873
rect -678 867 -620 873
rect -560 867 -502 873
rect -442 867 -384 873
rect -324 867 -266 873
rect -206 867 -148 873
rect -88 867 -30 873
rect 30 867 88 873
rect 148 867 206 873
rect 266 867 324 873
rect 384 867 442 873
rect 502 867 560 873
rect 620 867 678 873
rect 738 867 796 873
rect 856 867 914 873
rect 974 867 1032 873
rect 1092 867 1150 873
rect 1210 867 1268 873
rect 1328 867 1386 873
rect 1446 867 1504 873
rect 1564 867 1622 873
rect 1682 867 1740 873
rect 1800 867 1858 873
rect 1918 867 1976 873
rect 2036 867 2094 873
rect 2154 867 2212 873
rect 2272 867 2330 873
rect 2390 867 2448 873
rect 2508 867 2566 873
rect 2626 867 2684 873
rect 2744 867 2802 873
rect 2862 867 2920 873
rect -2920 799 -2862 805
rect -2802 799 -2744 805
rect -2684 799 -2626 805
rect -2566 799 -2508 805
rect -2448 799 -2390 805
rect -2330 799 -2272 805
rect -2212 799 -2154 805
rect -2094 799 -2036 805
rect -1976 799 -1918 805
rect -1858 799 -1800 805
rect -1740 799 -1682 805
rect -1622 799 -1564 805
rect -1504 799 -1446 805
rect -1386 799 -1328 805
rect -1268 799 -1210 805
rect -1150 799 -1092 805
rect -1032 799 -974 805
rect -914 799 -856 805
rect -796 799 -738 805
rect -678 799 -620 805
rect -560 799 -502 805
rect -442 799 -384 805
rect -324 799 -266 805
rect -206 799 -148 805
rect -88 799 -30 805
rect 30 799 88 805
rect 148 799 206 805
rect 266 799 324 805
rect 384 799 442 805
rect 502 799 560 805
rect 620 799 678 805
rect 738 799 796 805
rect 856 799 914 805
rect 974 799 1032 805
rect 1092 799 1150 805
rect 1210 799 1268 805
rect 1328 799 1386 805
rect 1446 799 1504 805
rect 1564 799 1622 805
rect 1682 799 1740 805
rect 1800 799 1858 805
rect 1918 799 1976 805
rect 2036 799 2094 805
rect 2154 799 2212 805
rect 2272 799 2330 805
rect 2390 799 2448 805
rect 2508 799 2566 805
rect 2626 799 2684 805
rect 2744 799 2802 805
rect 2862 799 2920 805
rect -2920 765 -2908 799
rect -2802 765 -2790 799
rect -2684 765 -2672 799
rect -2566 765 -2554 799
rect -2448 765 -2436 799
rect -2330 765 -2318 799
rect -2212 765 -2200 799
rect -2094 765 -2082 799
rect -1976 765 -1964 799
rect -1858 765 -1846 799
rect -1740 765 -1728 799
rect -1622 765 -1610 799
rect -1504 765 -1492 799
rect -1386 765 -1374 799
rect -1268 765 -1256 799
rect -1150 765 -1138 799
rect -1032 765 -1020 799
rect -914 765 -902 799
rect -796 765 -784 799
rect -678 765 -666 799
rect -560 765 -548 799
rect -442 765 -430 799
rect -324 765 -312 799
rect -206 765 -194 799
rect -88 765 -76 799
rect 30 765 42 799
rect 148 765 160 799
rect 266 765 278 799
rect 384 765 396 799
rect 502 765 514 799
rect 620 765 632 799
rect 738 765 750 799
rect 856 765 868 799
rect 974 765 986 799
rect 1092 765 1104 799
rect 1210 765 1222 799
rect 1328 765 1340 799
rect 1446 765 1458 799
rect 1564 765 1576 799
rect 1682 765 1694 799
rect 1800 765 1812 799
rect 1918 765 1930 799
rect 2036 765 2048 799
rect 2154 765 2166 799
rect 2272 765 2284 799
rect 2390 765 2402 799
rect 2508 765 2520 799
rect 2626 765 2638 799
rect 2744 765 2756 799
rect 2862 765 2874 799
rect -2920 759 -2862 765
rect -2802 759 -2744 765
rect -2684 759 -2626 765
rect -2566 759 -2508 765
rect -2448 759 -2390 765
rect -2330 759 -2272 765
rect -2212 759 -2154 765
rect -2094 759 -2036 765
rect -1976 759 -1918 765
rect -1858 759 -1800 765
rect -1740 759 -1682 765
rect -1622 759 -1564 765
rect -1504 759 -1446 765
rect -1386 759 -1328 765
rect -1268 759 -1210 765
rect -1150 759 -1092 765
rect -1032 759 -974 765
rect -914 759 -856 765
rect -796 759 -738 765
rect -678 759 -620 765
rect -560 759 -502 765
rect -442 759 -384 765
rect -324 759 -266 765
rect -206 759 -148 765
rect -88 759 -30 765
rect 30 759 88 765
rect 148 759 206 765
rect 266 759 324 765
rect 384 759 442 765
rect 502 759 560 765
rect 620 759 678 765
rect 738 759 796 765
rect 856 759 914 765
rect 974 759 1032 765
rect 1092 759 1150 765
rect 1210 759 1268 765
rect 1328 759 1386 765
rect 1446 759 1504 765
rect 1564 759 1622 765
rect 1682 759 1740 765
rect 1800 759 1858 765
rect 1918 759 1976 765
rect 2036 759 2094 765
rect 2154 759 2212 765
rect 2272 759 2330 765
rect 2390 759 2448 765
rect 2508 759 2566 765
rect 2626 759 2684 765
rect 2744 759 2802 765
rect 2862 759 2920 765
rect -2920 71 -2862 77
rect -2802 71 -2744 77
rect -2684 71 -2626 77
rect -2566 71 -2508 77
rect -2448 71 -2390 77
rect -2330 71 -2272 77
rect -2212 71 -2154 77
rect -2094 71 -2036 77
rect -1976 71 -1918 77
rect -1858 71 -1800 77
rect -1740 71 -1682 77
rect -1622 71 -1564 77
rect -1504 71 -1446 77
rect -1386 71 -1328 77
rect -1268 71 -1210 77
rect -1150 71 -1092 77
rect -1032 71 -974 77
rect -914 71 -856 77
rect -796 71 -738 77
rect -678 71 -620 77
rect -560 71 -502 77
rect -442 71 -384 77
rect -324 71 -266 77
rect -206 71 -148 77
rect -88 71 -30 77
rect 30 71 88 77
rect 148 71 206 77
rect 266 71 324 77
rect 384 71 442 77
rect 502 71 560 77
rect 620 71 678 77
rect 738 71 796 77
rect 856 71 914 77
rect 974 71 1032 77
rect 1092 71 1150 77
rect 1210 71 1268 77
rect 1328 71 1386 77
rect 1446 71 1504 77
rect 1564 71 1622 77
rect 1682 71 1740 77
rect 1800 71 1858 77
rect 1918 71 1976 77
rect 2036 71 2094 77
rect 2154 71 2212 77
rect 2272 71 2330 77
rect 2390 71 2448 77
rect 2508 71 2566 77
rect 2626 71 2684 77
rect 2744 71 2802 77
rect 2862 71 2920 77
rect -2920 37 -2908 71
rect -2802 37 -2790 71
rect -2684 37 -2672 71
rect -2566 37 -2554 71
rect -2448 37 -2436 71
rect -2330 37 -2318 71
rect -2212 37 -2200 71
rect -2094 37 -2082 71
rect -1976 37 -1964 71
rect -1858 37 -1846 71
rect -1740 37 -1728 71
rect -1622 37 -1610 71
rect -1504 37 -1492 71
rect -1386 37 -1374 71
rect -1268 37 -1256 71
rect -1150 37 -1138 71
rect -1032 37 -1020 71
rect -914 37 -902 71
rect -796 37 -784 71
rect -678 37 -666 71
rect -560 37 -548 71
rect -442 37 -430 71
rect -324 37 -312 71
rect -206 37 -194 71
rect -88 37 -76 71
rect 30 37 42 71
rect 148 37 160 71
rect 266 37 278 71
rect 384 37 396 71
rect 502 37 514 71
rect 620 37 632 71
rect 738 37 750 71
rect 856 37 868 71
rect 974 37 986 71
rect 1092 37 1104 71
rect 1210 37 1222 71
rect 1328 37 1340 71
rect 1446 37 1458 71
rect 1564 37 1576 71
rect 1682 37 1694 71
rect 1800 37 1812 71
rect 1918 37 1930 71
rect 2036 37 2048 71
rect 2154 37 2166 71
rect 2272 37 2284 71
rect 2390 37 2402 71
rect 2508 37 2520 71
rect 2626 37 2638 71
rect 2744 37 2756 71
rect 2862 37 2874 71
rect -2920 31 -2862 37
rect -2802 31 -2744 37
rect -2684 31 -2626 37
rect -2566 31 -2508 37
rect -2448 31 -2390 37
rect -2330 31 -2272 37
rect -2212 31 -2154 37
rect -2094 31 -2036 37
rect -1976 31 -1918 37
rect -1858 31 -1800 37
rect -1740 31 -1682 37
rect -1622 31 -1564 37
rect -1504 31 -1446 37
rect -1386 31 -1328 37
rect -1268 31 -1210 37
rect -1150 31 -1092 37
rect -1032 31 -974 37
rect -914 31 -856 37
rect -796 31 -738 37
rect -678 31 -620 37
rect -560 31 -502 37
rect -442 31 -384 37
rect -324 31 -266 37
rect -206 31 -148 37
rect -88 31 -30 37
rect 30 31 88 37
rect 148 31 206 37
rect 266 31 324 37
rect 384 31 442 37
rect 502 31 560 37
rect 620 31 678 37
rect 738 31 796 37
rect 856 31 914 37
rect 974 31 1032 37
rect 1092 31 1150 37
rect 1210 31 1268 37
rect 1328 31 1386 37
rect 1446 31 1504 37
rect 1564 31 1622 37
rect 1682 31 1740 37
rect 1800 31 1858 37
rect 1918 31 1976 37
rect 2036 31 2094 37
rect 2154 31 2212 37
rect 2272 31 2330 37
rect 2390 31 2448 37
rect 2508 31 2566 37
rect 2626 31 2684 37
rect 2744 31 2802 37
rect 2862 31 2920 37
rect -2920 -37 -2862 -31
rect -2802 -37 -2744 -31
rect -2684 -37 -2626 -31
rect -2566 -37 -2508 -31
rect -2448 -37 -2390 -31
rect -2330 -37 -2272 -31
rect -2212 -37 -2154 -31
rect -2094 -37 -2036 -31
rect -1976 -37 -1918 -31
rect -1858 -37 -1800 -31
rect -1740 -37 -1682 -31
rect -1622 -37 -1564 -31
rect -1504 -37 -1446 -31
rect -1386 -37 -1328 -31
rect -1268 -37 -1210 -31
rect -1150 -37 -1092 -31
rect -1032 -37 -974 -31
rect -914 -37 -856 -31
rect -796 -37 -738 -31
rect -678 -37 -620 -31
rect -560 -37 -502 -31
rect -442 -37 -384 -31
rect -324 -37 -266 -31
rect -206 -37 -148 -31
rect -88 -37 -30 -31
rect 30 -37 88 -31
rect 148 -37 206 -31
rect 266 -37 324 -31
rect 384 -37 442 -31
rect 502 -37 560 -31
rect 620 -37 678 -31
rect 738 -37 796 -31
rect 856 -37 914 -31
rect 974 -37 1032 -31
rect 1092 -37 1150 -31
rect 1210 -37 1268 -31
rect 1328 -37 1386 -31
rect 1446 -37 1504 -31
rect 1564 -37 1622 -31
rect 1682 -37 1740 -31
rect 1800 -37 1858 -31
rect 1918 -37 1976 -31
rect 2036 -37 2094 -31
rect 2154 -37 2212 -31
rect 2272 -37 2330 -31
rect 2390 -37 2448 -31
rect 2508 -37 2566 -31
rect 2626 -37 2684 -31
rect 2744 -37 2802 -31
rect 2862 -37 2920 -31
rect -2920 -71 -2908 -37
rect -2802 -71 -2790 -37
rect -2684 -71 -2672 -37
rect -2566 -71 -2554 -37
rect -2448 -71 -2436 -37
rect -2330 -71 -2318 -37
rect -2212 -71 -2200 -37
rect -2094 -71 -2082 -37
rect -1976 -71 -1964 -37
rect -1858 -71 -1846 -37
rect -1740 -71 -1728 -37
rect -1622 -71 -1610 -37
rect -1504 -71 -1492 -37
rect -1386 -71 -1374 -37
rect -1268 -71 -1256 -37
rect -1150 -71 -1138 -37
rect -1032 -71 -1020 -37
rect -914 -71 -902 -37
rect -796 -71 -784 -37
rect -678 -71 -666 -37
rect -560 -71 -548 -37
rect -442 -71 -430 -37
rect -324 -71 -312 -37
rect -206 -71 -194 -37
rect -88 -71 -76 -37
rect 30 -71 42 -37
rect 148 -71 160 -37
rect 266 -71 278 -37
rect 384 -71 396 -37
rect 502 -71 514 -37
rect 620 -71 632 -37
rect 738 -71 750 -37
rect 856 -71 868 -37
rect 974 -71 986 -37
rect 1092 -71 1104 -37
rect 1210 -71 1222 -37
rect 1328 -71 1340 -37
rect 1446 -71 1458 -37
rect 1564 -71 1576 -37
rect 1682 -71 1694 -37
rect 1800 -71 1812 -37
rect 1918 -71 1930 -37
rect 2036 -71 2048 -37
rect 2154 -71 2166 -37
rect 2272 -71 2284 -37
rect 2390 -71 2402 -37
rect 2508 -71 2520 -37
rect 2626 -71 2638 -37
rect 2744 -71 2756 -37
rect 2862 -71 2874 -37
rect -2920 -77 -2862 -71
rect -2802 -77 -2744 -71
rect -2684 -77 -2626 -71
rect -2566 -77 -2508 -71
rect -2448 -77 -2390 -71
rect -2330 -77 -2272 -71
rect -2212 -77 -2154 -71
rect -2094 -77 -2036 -71
rect -1976 -77 -1918 -71
rect -1858 -77 -1800 -71
rect -1740 -77 -1682 -71
rect -1622 -77 -1564 -71
rect -1504 -77 -1446 -71
rect -1386 -77 -1328 -71
rect -1268 -77 -1210 -71
rect -1150 -77 -1092 -71
rect -1032 -77 -974 -71
rect -914 -77 -856 -71
rect -796 -77 -738 -71
rect -678 -77 -620 -71
rect -560 -77 -502 -71
rect -442 -77 -384 -71
rect -324 -77 -266 -71
rect -206 -77 -148 -71
rect -88 -77 -30 -71
rect 30 -77 88 -71
rect 148 -77 206 -71
rect 266 -77 324 -71
rect 384 -77 442 -71
rect 502 -77 560 -71
rect 620 -77 678 -71
rect 738 -77 796 -71
rect 856 -77 914 -71
rect 974 -77 1032 -71
rect 1092 -77 1150 -71
rect 1210 -77 1268 -71
rect 1328 -77 1386 -71
rect 1446 -77 1504 -71
rect 1564 -77 1622 -71
rect 1682 -77 1740 -71
rect 1800 -77 1858 -71
rect 1918 -77 1976 -71
rect 2036 -77 2094 -71
rect 2154 -77 2212 -71
rect 2272 -77 2330 -71
rect 2390 -77 2448 -71
rect 2508 -77 2566 -71
rect 2626 -77 2684 -71
rect 2744 -77 2802 -71
rect 2862 -77 2920 -71
rect -2920 -765 -2862 -759
rect -2802 -765 -2744 -759
rect -2684 -765 -2626 -759
rect -2566 -765 -2508 -759
rect -2448 -765 -2390 -759
rect -2330 -765 -2272 -759
rect -2212 -765 -2154 -759
rect -2094 -765 -2036 -759
rect -1976 -765 -1918 -759
rect -1858 -765 -1800 -759
rect -1740 -765 -1682 -759
rect -1622 -765 -1564 -759
rect -1504 -765 -1446 -759
rect -1386 -765 -1328 -759
rect -1268 -765 -1210 -759
rect -1150 -765 -1092 -759
rect -1032 -765 -974 -759
rect -914 -765 -856 -759
rect -796 -765 -738 -759
rect -678 -765 -620 -759
rect -560 -765 -502 -759
rect -442 -765 -384 -759
rect -324 -765 -266 -759
rect -206 -765 -148 -759
rect -88 -765 -30 -759
rect 30 -765 88 -759
rect 148 -765 206 -759
rect 266 -765 324 -759
rect 384 -765 442 -759
rect 502 -765 560 -759
rect 620 -765 678 -759
rect 738 -765 796 -759
rect 856 -765 914 -759
rect 974 -765 1032 -759
rect 1092 -765 1150 -759
rect 1210 -765 1268 -759
rect 1328 -765 1386 -759
rect 1446 -765 1504 -759
rect 1564 -765 1622 -759
rect 1682 -765 1740 -759
rect 1800 -765 1858 -759
rect 1918 -765 1976 -759
rect 2036 -765 2094 -759
rect 2154 -765 2212 -759
rect 2272 -765 2330 -759
rect 2390 -765 2448 -759
rect 2508 -765 2566 -759
rect 2626 -765 2684 -759
rect 2744 -765 2802 -759
rect 2862 -765 2920 -759
rect -2920 -799 -2908 -765
rect -2802 -799 -2790 -765
rect -2684 -799 -2672 -765
rect -2566 -799 -2554 -765
rect -2448 -799 -2436 -765
rect -2330 -799 -2318 -765
rect -2212 -799 -2200 -765
rect -2094 -799 -2082 -765
rect -1976 -799 -1964 -765
rect -1858 -799 -1846 -765
rect -1740 -799 -1728 -765
rect -1622 -799 -1610 -765
rect -1504 -799 -1492 -765
rect -1386 -799 -1374 -765
rect -1268 -799 -1256 -765
rect -1150 -799 -1138 -765
rect -1032 -799 -1020 -765
rect -914 -799 -902 -765
rect -796 -799 -784 -765
rect -678 -799 -666 -765
rect -560 -799 -548 -765
rect -442 -799 -430 -765
rect -324 -799 -312 -765
rect -206 -799 -194 -765
rect -88 -799 -76 -765
rect 30 -799 42 -765
rect 148 -799 160 -765
rect 266 -799 278 -765
rect 384 -799 396 -765
rect 502 -799 514 -765
rect 620 -799 632 -765
rect 738 -799 750 -765
rect 856 -799 868 -765
rect 974 -799 986 -765
rect 1092 -799 1104 -765
rect 1210 -799 1222 -765
rect 1328 -799 1340 -765
rect 1446 -799 1458 -765
rect 1564 -799 1576 -765
rect 1682 -799 1694 -765
rect 1800 -799 1812 -765
rect 1918 -799 1930 -765
rect 2036 -799 2048 -765
rect 2154 -799 2166 -765
rect 2272 -799 2284 -765
rect 2390 -799 2402 -765
rect 2508 -799 2520 -765
rect 2626 -799 2638 -765
rect 2744 -799 2756 -765
rect 2862 -799 2874 -765
rect -2920 -805 -2862 -799
rect -2802 -805 -2744 -799
rect -2684 -805 -2626 -799
rect -2566 -805 -2508 -799
rect -2448 -805 -2390 -799
rect -2330 -805 -2272 -799
rect -2212 -805 -2154 -799
rect -2094 -805 -2036 -799
rect -1976 -805 -1918 -799
rect -1858 -805 -1800 -799
rect -1740 -805 -1682 -799
rect -1622 -805 -1564 -799
rect -1504 -805 -1446 -799
rect -1386 -805 -1328 -799
rect -1268 -805 -1210 -799
rect -1150 -805 -1092 -799
rect -1032 -805 -974 -799
rect -914 -805 -856 -799
rect -796 -805 -738 -799
rect -678 -805 -620 -799
rect -560 -805 -502 -799
rect -442 -805 -384 -799
rect -324 -805 -266 -799
rect -206 -805 -148 -799
rect -88 -805 -30 -799
rect 30 -805 88 -799
rect 148 -805 206 -799
rect 266 -805 324 -799
rect 384 -805 442 -799
rect 502 -805 560 -799
rect 620 -805 678 -799
rect 738 -805 796 -799
rect 856 -805 914 -799
rect 974 -805 1032 -799
rect 1092 -805 1150 -799
rect 1210 -805 1268 -799
rect 1328 -805 1386 -799
rect 1446 -805 1504 -799
rect 1564 -805 1622 -799
rect 1682 -805 1740 -799
rect 1800 -805 1858 -799
rect 1918 -805 1976 -799
rect 2036 -805 2094 -799
rect 2154 -805 2212 -799
rect 2272 -805 2330 -799
rect 2390 -805 2448 -799
rect 2508 -805 2566 -799
rect 2626 -805 2684 -799
rect 2744 -805 2802 -799
rect 2862 -805 2920 -799
rect -2920 -873 -2862 -867
rect -2802 -873 -2744 -867
rect -2684 -873 -2626 -867
rect -2566 -873 -2508 -867
rect -2448 -873 -2390 -867
rect -2330 -873 -2272 -867
rect -2212 -873 -2154 -867
rect -2094 -873 -2036 -867
rect -1976 -873 -1918 -867
rect -1858 -873 -1800 -867
rect -1740 -873 -1682 -867
rect -1622 -873 -1564 -867
rect -1504 -873 -1446 -867
rect -1386 -873 -1328 -867
rect -1268 -873 -1210 -867
rect -1150 -873 -1092 -867
rect -1032 -873 -974 -867
rect -914 -873 -856 -867
rect -796 -873 -738 -867
rect -678 -873 -620 -867
rect -560 -873 -502 -867
rect -442 -873 -384 -867
rect -324 -873 -266 -867
rect -206 -873 -148 -867
rect -88 -873 -30 -867
rect 30 -873 88 -867
rect 148 -873 206 -867
rect 266 -873 324 -867
rect 384 -873 442 -867
rect 502 -873 560 -867
rect 620 -873 678 -867
rect 738 -873 796 -867
rect 856 -873 914 -867
rect 974 -873 1032 -867
rect 1092 -873 1150 -867
rect 1210 -873 1268 -867
rect 1328 -873 1386 -867
rect 1446 -873 1504 -867
rect 1564 -873 1622 -867
rect 1682 -873 1740 -867
rect 1800 -873 1858 -867
rect 1918 -873 1976 -867
rect 2036 -873 2094 -867
rect 2154 -873 2212 -867
rect 2272 -873 2330 -867
rect 2390 -873 2448 -867
rect 2508 -873 2566 -867
rect 2626 -873 2684 -867
rect 2744 -873 2802 -867
rect 2862 -873 2920 -867
rect -2920 -907 -2908 -873
rect -2802 -907 -2790 -873
rect -2684 -907 -2672 -873
rect -2566 -907 -2554 -873
rect -2448 -907 -2436 -873
rect -2330 -907 -2318 -873
rect -2212 -907 -2200 -873
rect -2094 -907 -2082 -873
rect -1976 -907 -1964 -873
rect -1858 -907 -1846 -873
rect -1740 -907 -1728 -873
rect -1622 -907 -1610 -873
rect -1504 -907 -1492 -873
rect -1386 -907 -1374 -873
rect -1268 -907 -1256 -873
rect -1150 -907 -1138 -873
rect -1032 -907 -1020 -873
rect -914 -907 -902 -873
rect -796 -907 -784 -873
rect -678 -907 -666 -873
rect -560 -907 -548 -873
rect -442 -907 -430 -873
rect -324 -907 -312 -873
rect -206 -907 -194 -873
rect -88 -907 -76 -873
rect 30 -907 42 -873
rect 148 -907 160 -873
rect 266 -907 278 -873
rect 384 -907 396 -873
rect 502 -907 514 -873
rect 620 -907 632 -873
rect 738 -907 750 -873
rect 856 -907 868 -873
rect 974 -907 986 -873
rect 1092 -907 1104 -873
rect 1210 -907 1222 -873
rect 1328 -907 1340 -873
rect 1446 -907 1458 -873
rect 1564 -907 1576 -873
rect 1682 -907 1694 -873
rect 1800 -907 1812 -873
rect 1918 -907 1930 -873
rect 2036 -907 2048 -873
rect 2154 -907 2166 -873
rect 2272 -907 2284 -873
rect 2390 -907 2402 -873
rect 2508 -907 2520 -873
rect 2626 -907 2638 -873
rect 2744 -907 2756 -873
rect 2862 -907 2874 -873
rect -2920 -913 -2862 -907
rect -2802 -913 -2744 -907
rect -2684 -913 -2626 -907
rect -2566 -913 -2508 -907
rect -2448 -913 -2390 -907
rect -2330 -913 -2272 -907
rect -2212 -913 -2154 -907
rect -2094 -913 -2036 -907
rect -1976 -913 -1918 -907
rect -1858 -913 -1800 -907
rect -1740 -913 -1682 -907
rect -1622 -913 -1564 -907
rect -1504 -913 -1446 -907
rect -1386 -913 -1328 -907
rect -1268 -913 -1210 -907
rect -1150 -913 -1092 -907
rect -1032 -913 -974 -907
rect -914 -913 -856 -907
rect -796 -913 -738 -907
rect -678 -913 -620 -907
rect -560 -913 -502 -907
rect -442 -913 -384 -907
rect -324 -913 -266 -907
rect -206 -913 -148 -907
rect -88 -913 -30 -907
rect 30 -913 88 -907
rect 148 -913 206 -907
rect 266 -913 324 -907
rect 384 -913 442 -907
rect 502 -913 560 -907
rect 620 -913 678 -907
rect 738 -913 796 -907
rect 856 -913 914 -907
rect 974 -913 1032 -907
rect 1092 -913 1150 -907
rect 1210 -913 1268 -907
rect 1328 -913 1386 -907
rect 1446 -913 1504 -907
rect 1564 -913 1622 -907
rect 1682 -913 1740 -907
rect 1800 -913 1858 -907
rect 1918 -913 1976 -907
rect 2036 -913 2094 -907
rect 2154 -913 2212 -907
rect 2272 -913 2330 -907
rect 2390 -913 2448 -907
rect 2508 -913 2566 -907
rect 2626 -913 2684 -907
rect 2744 -913 2802 -907
rect 2862 -913 2920 -907
rect -2920 -1601 -2862 -1595
rect -2802 -1601 -2744 -1595
rect -2684 -1601 -2626 -1595
rect -2566 -1601 -2508 -1595
rect -2448 -1601 -2390 -1595
rect -2330 -1601 -2272 -1595
rect -2212 -1601 -2154 -1595
rect -2094 -1601 -2036 -1595
rect -1976 -1601 -1918 -1595
rect -1858 -1601 -1800 -1595
rect -1740 -1601 -1682 -1595
rect -1622 -1601 -1564 -1595
rect -1504 -1601 -1446 -1595
rect -1386 -1601 -1328 -1595
rect -1268 -1601 -1210 -1595
rect -1150 -1601 -1092 -1595
rect -1032 -1601 -974 -1595
rect -914 -1601 -856 -1595
rect -796 -1601 -738 -1595
rect -678 -1601 -620 -1595
rect -560 -1601 -502 -1595
rect -442 -1601 -384 -1595
rect -324 -1601 -266 -1595
rect -206 -1601 -148 -1595
rect -88 -1601 -30 -1595
rect 30 -1601 88 -1595
rect 148 -1601 206 -1595
rect 266 -1601 324 -1595
rect 384 -1601 442 -1595
rect 502 -1601 560 -1595
rect 620 -1601 678 -1595
rect 738 -1601 796 -1595
rect 856 -1601 914 -1595
rect 974 -1601 1032 -1595
rect 1092 -1601 1150 -1595
rect 1210 -1601 1268 -1595
rect 1328 -1601 1386 -1595
rect 1446 -1601 1504 -1595
rect 1564 -1601 1622 -1595
rect 1682 -1601 1740 -1595
rect 1800 -1601 1858 -1595
rect 1918 -1601 1976 -1595
rect 2036 -1601 2094 -1595
rect 2154 -1601 2212 -1595
rect 2272 -1601 2330 -1595
rect 2390 -1601 2448 -1595
rect 2508 -1601 2566 -1595
rect 2626 -1601 2684 -1595
rect 2744 -1601 2802 -1595
rect 2862 -1601 2920 -1595
rect -2920 -1635 -2908 -1601
rect -2802 -1635 -2790 -1601
rect -2684 -1635 -2672 -1601
rect -2566 -1635 -2554 -1601
rect -2448 -1635 -2436 -1601
rect -2330 -1635 -2318 -1601
rect -2212 -1635 -2200 -1601
rect -2094 -1635 -2082 -1601
rect -1976 -1635 -1964 -1601
rect -1858 -1635 -1846 -1601
rect -1740 -1635 -1728 -1601
rect -1622 -1635 -1610 -1601
rect -1504 -1635 -1492 -1601
rect -1386 -1635 -1374 -1601
rect -1268 -1635 -1256 -1601
rect -1150 -1635 -1138 -1601
rect -1032 -1635 -1020 -1601
rect -914 -1635 -902 -1601
rect -796 -1635 -784 -1601
rect -678 -1635 -666 -1601
rect -560 -1635 -548 -1601
rect -442 -1635 -430 -1601
rect -324 -1635 -312 -1601
rect -206 -1635 -194 -1601
rect -88 -1635 -76 -1601
rect 30 -1635 42 -1601
rect 148 -1635 160 -1601
rect 266 -1635 278 -1601
rect 384 -1635 396 -1601
rect 502 -1635 514 -1601
rect 620 -1635 632 -1601
rect 738 -1635 750 -1601
rect 856 -1635 868 -1601
rect 974 -1635 986 -1601
rect 1092 -1635 1104 -1601
rect 1210 -1635 1222 -1601
rect 1328 -1635 1340 -1601
rect 1446 -1635 1458 -1601
rect 1564 -1635 1576 -1601
rect 1682 -1635 1694 -1601
rect 1800 -1635 1812 -1601
rect 1918 -1635 1930 -1601
rect 2036 -1635 2048 -1601
rect 2154 -1635 2166 -1601
rect 2272 -1635 2284 -1601
rect 2390 -1635 2402 -1601
rect 2508 -1635 2520 -1601
rect 2626 -1635 2638 -1601
rect 2744 -1635 2756 -1601
rect 2862 -1635 2874 -1601
rect -2920 -1641 -2862 -1635
rect -2802 -1641 -2744 -1635
rect -2684 -1641 -2626 -1635
rect -2566 -1641 -2508 -1635
rect -2448 -1641 -2390 -1635
rect -2330 -1641 -2272 -1635
rect -2212 -1641 -2154 -1635
rect -2094 -1641 -2036 -1635
rect -1976 -1641 -1918 -1635
rect -1858 -1641 -1800 -1635
rect -1740 -1641 -1682 -1635
rect -1622 -1641 -1564 -1635
rect -1504 -1641 -1446 -1635
rect -1386 -1641 -1328 -1635
rect -1268 -1641 -1210 -1635
rect -1150 -1641 -1092 -1635
rect -1032 -1641 -974 -1635
rect -914 -1641 -856 -1635
rect -796 -1641 -738 -1635
rect -678 -1641 -620 -1635
rect -560 -1641 -502 -1635
rect -442 -1641 -384 -1635
rect -324 -1641 -266 -1635
rect -206 -1641 -148 -1635
rect -88 -1641 -30 -1635
rect 30 -1641 88 -1635
rect 148 -1641 206 -1635
rect 266 -1641 324 -1635
rect 384 -1641 442 -1635
rect 502 -1641 560 -1635
rect 620 -1641 678 -1635
rect 738 -1641 796 -1635
rect 856 -1641 914 -1635
rect 974 -1641 1032 -1635
rect 1092 -1641 1150 -1635
rect 1210 -1641 1268 -1635
rect 1328 -1641 1386 -1635
rect 1446 -1641 1504 -1635
rect 1564 -1641 1622 -1635
rect 1682 -1641 1740 -1635
rect 1800 -1641 1858 -1635
rect 1918 -1641 1976 -1635
rect 2036 -1641 2094 -1635
rect 2154 -1641 2212 -1635
rect 2272 -1641 2330 -1635
rect 2390 -1641 2448 -1635
rect 2508 -1641 2566 -1635
rect 2626 -1641 2684 -1635
rect 2744 -1641 2802 -1635
rect 2862 -1641 2920 -1635
<< nwell >>
rect -3117 -1773 3117 1773
<< pmos >>
rect -2921 954 -2861 1554
rect -2803 954 -2743 1554
rect -2685 954 -2625 1554
rect -2567 954 -2507 1554
rect -2449 954 -2389 1554
rect -2331 954 -2271 1554
rect -2213 954 -2153 1554
rect -2095 954 -2035 1554
rect -1977 954 -1917 1554
rect -1859 954 -1799 1554
rect -1741 954 -1681 1554
rect -1623 954 -1563 1554
rect -1505 954 -1445 1554
rect -1387 954 -1327 1554
rect -1269 954 -1209 1554
rect -1151 954 -1091 1554
rect -1033 954 -973 1554
rect -915 954 -855 1554
rect -797 954 -737 1554
rect -679 954 -619 1554
rect -561 954 -501 1554
rect -443 954 -383 1554
rect -325 954 -265 1554
rect -207 954 -147 1554
rect -89 954 -29 1554
rect 29 954 89 1554
rect 147 954 207 1554
rect 265 954 325 1554
rect 383 954 443 1554
rect 501 954 561 1554
rect 619 954 679 1554
rect 737 954 797 1554
rect 855 954 915 1554
rect 973 954 1033 1554
rect 1091 954 1151 1554
rect 1209 954 1269 1554
rect 1327 954 1387 1554
rect 1445 954 1505 1554
rect 1563 954 1623 1554
rect 1681 954 1741 1554
rect 1799 954 1859 1554
rect 1917 954 1977 1554
rect 2035 954 2095 1554
rect 2153 954 2213 1554
rect 2271 954 2331 1554
rect 2389 954 2449 1554
rect 2507 954 2567 1554
rect 2625 954 2685 1554
rect 2743 954 2803 1554
rect 2861 954 2921 1554
rect -2921 118 -2861 718
rect -2803 118 -2743 718
rect -2685 118 -2625 718
rect -2567 118 -2507 718
rect -2449 118 -2389 718
rect -2331 118 -2271 718
rect -2213 118 -2153 718
rect -2095 118 -2035 718
rect -1977 118 -1917 718
rect -1859 118 -1799 718
rect -1741 118 -1681 718
rect -1623 118 -1563 718
rect -1505 118 -1445 718
rect -1387 118 -1327 718
rect -1269 118 -1209 718
rect -1151 118 -1091 718
rect -1033 118 -973 718
rect -915 118 -855 718
rect -797 118 -737 718
rect -679 118 -619 718
rect -561 118 -501 718
rect -443 118 -383 718
rect -325 118 -265 718
rect -207 118 -147 718
rect -89 118 -29 718
rect 29 118 89 718
rect 147 118 207 718
rect 265 118 325 718
rect 383 118 443 718
rect 501 118 561 718
rect 619 118 679 718
rect 737 118 797 718
rect 855 118 915 718
rect 973 118 1033 718
rect 1091 118 1151 718
rect 1209 118 1269 718
rect 1327 118 1387 718
rect 1445 118 1505 718
rect 1563 118 1623 718
rect 1681 118 1741 718
rect 1799 118 1859 718
rect 1917 118 1977 718
rect 2035 118 2095 718
rect 2153 118 2213 718
rect 2271 118 2331 718
rect 2389 118 2449 718
rect 2507 118 2567 718
rect 2625 118 2685 718
rect 2743 118 2803 718
rect 2861 118 2921 718
rect -2921 -718 -2861 -118
rect -2803 -718 -2743 -118
rect -2685 -718 -2625 -118
rect -2567 -718 -2507 -118
rect -2449 -718 -2389 -118
rect -2331 -718 -2271 -118
rect -2213 -718 -2153 -118
rect -2095 -718 -2035 -118
rect -1977 -718 -1917 -118
rect -1859 -718 -1799 -118
rect -1741 -718 -1681 -118
rect -1623 -718 -1563 -118
rect -1505 -718 -1445 -118
rect -1387 -718 -1327 -118
rect -1269 -718 -1209 -118
rect -1151 -718 -1091 -118
rect -1033 -718 -973 -118
rect -915 -718 -855 -118
rect -797 -718 -737 -118
rect -679 -718 -619 -118
rect -561 -718 -501 -118
rect -443 -718 -383 -118
rect -325 -718 -265 -118
rect -207 -718 -147 -118
rect -89 -718 -29 -118
rect 29 -718 89 -118
rect 147 -718 207 -118
rect 265 -718 325 -118
rect 383 -718 443 -118
rect 501 -718 561 -118
rect 619 -718 679 -118
rect 737 -718 797 -118
rect 855 -718 915 -118
rect 973 -718 1033 -118
rect 1091 -718 1151 -118
rect 1209 -718 1269 -118
rect 1327 -718 1387 -118
rect 1445 -718 1505 -118
rect 1563 -718 1623 -118
rect 1681 -718 1741 -118
rect 1799 -718 1859 -118
rect 1917 -718 1977 -118
rect 2035 -718 2095 -118
rect 2153 -718 2213 -118
rect 2271 -718 2331 -118
rect 2389 -718 2449 -118
rect 2507 -718 2567 -118
rect 2625 -718 2685 -118
rect 2743 -718 2803 -118
rect 2861 -718 2921 -118
rect -2921 -1554 -2861 -954
rect -2803 -1554 -2743 -954
rect -2685 -1554 -2625 -954
rect -2567 -1554 -2507 -954
rect -2449 -1554 -2389 -954
rect -2331 -1554 -2271 -954
rect -2213 -1554 -2153 -954
rect -2095 -1554 -2035 -954
rect -1977 -1554 -1917 -954
rect -1859 -1554 -1799 -954
rect -1741 -1554 -1681 -954
rect -1623 -1554 -1563 -954
rect -1505 -1554 -1445 -954
rect -1387 -1554 -1327 -954
rect -1269 -1554 -1209 -954
rect -1151 -1554 -1091 -954
rect -1033 -1554 -973 -954
rect -915 -1554 -855 -954
rect -797 -1554 -737 -954
rect -679 -1554 -619 -954
rect -561 -1554 -501 -954
rect -443 -1554 -383 -954
rect -325 -1554 -265 -954
rect -207 -1554 -147 -954
rect -89 -1554 -29 -954
rect 29 -1554 89 -954
rect 147 -1554 207 -954
rect 265 -1554 325 -954
rect 383 -1554 443 -954
rect 501 -1554 561 -954
rect 619 -1554 679 -954
rect 737 -1554 797 -954
rect 855 -1554 915 -954
rect 973 -1554 1033 -954
rect 1091 -1554 1151 -954
rect 1209 -1554 1269 -954
rect 1327 -1554 1387 -954
rect 1445 -1554 1505 -954
rect 1563 -1554 1623 -954
rect 1681 -1554 1741 -954
rect 1799 -1554 1859 -954
rect 1917 -1554 1977 -954
rect 2035 -1554 2095 -954
rect 2153 -1554 2213 -954
rect 2271 -1554 2331 -954
rect 2389 -1554 2449 -954
rect 2507 -1554 2567 -954
rect 2625 -1554 2685 -954
rect 2743 -1554 2803 -954
rect 2861 -1554 2921 -954
<< pdiff >>
rect -2979 1542 -2921 1554
rect -2979 966 -2967 1542
rect -2933 966 -2921 1542
rect -2979 954 -2921 966
rect -2861 1542 -2803 1554
rect -2861 966 -2849 1542
rect -2815 966 -2803 1542
rect -2861 954 -2803 966
rect -2743 1542 -2685 1554
rect -2743 966 -2731 1542
rect -2697 966 -2685 1542
rect -2743 954 -2685 966
rect -2625 1542 -2567 1554
rect -2625 966 -2613 1542
rect -2579 966 -2567 1542
rect -2625 954 -2567 966
rect -2507 1542 -2449 1554
rect -2507 966 -2495 1542
rect -2461 966 -2449 1542
rect -2507 954 -2449 966
rect -2389 1542 -2331 1554
rect -2389 966 -2377 1542
rect -2343 966 -2331 1542
rect -2389 954 -2331 966
rect -2271 1542 -2213 1554
rect -2271 966 -2259 1542
rect -2225 966 -2213 1542
rect -2271 954 -2213 966
rect -2153 1542 -2095 1554
rect -2153 966 -2141 1542
rect -2107 966 -2095 1542
rect -2153 954 -2095 966
rect -2035 1542 -1977 1554
rect -2035 966 -2023 1542
rect -1989 966 -1977 1542
rect -2035 954 -1977 966
rect -1917 1542 -1859 1554
rect -1917 966 -1905 1542
rect -1871 966 -1859 1542
rect -1917 954 -1859 966
rect -1799 1542 -1741 1554
rect -1799 966 -1787 1542
rect -1753 966 -1741 1542
rect -1799 954 -1741 966
rect -1681 1542 -1623 1554
rect -1681 966 -1669 1542
rect -1635 966 -1623 1542
rect -1681 954 -1623 966
rect -1563 1542 -1505 1554
rect -1563 966 -1551 1542
rect -1517 966 -1505 1542
rect -1563 954 -1505 966
rect -1445 1542 -1387 1554
rect -1445 966 -1433 1542
rect -1399 966 -1387 1542
rect -1445 954 -1387 966
rect -1327 1542 -1269 1554
rect -1327 966 -1315 1542
rect -1281 966 -1269 1542
rect -1327 954 -1269 966
rect -1209 1542 -1151 1554
rect -1209 966 -1197 1542
rect -1163 966 -1151 1542
rect -1209 954 -1151 966
rect -1091 1542 -1033 1554
rect -1091 966 -1079 1542
rect -1045 966 -1033 1542
rect -1091 954 -1033 966
rect -973 1542 -915 1554
rect -973 966 -961 1542
rect -927 966 -915 1542
rect -973 954 -915 966
rect -855 1542 -797 1554
rect -855 966 -843 1542
rect -809 966 -797 1542
rect -855 954 -797 966
rect -737 1542 -679 1554
rect -737 966 -725 1542
rect -691 966 -679 1542
rect -737 954 -679 966
rect -619 1542 -561 1554
rect -619 966 -607 1542
rect -573 966 -561 1542
rect -619 954 -561 966
rect -501 1542 -443 1554
rect -501 966 -489 1542
rect -455 966 -443 1542
rect -501 954 -443 966
rect -383 1542 -325 1554
rect -383 966 -371 1542
rect -337 966 -325 1542
rect -383 954 -325 966
rect -265 1542 -207 1554
rect -265 966 -253 1542
rect -219 966 -207 1542
rect -265 954 -207 966
rect -147 1542 -89 1554
rect -147 966 -135 1542
rect -101 966 -89 1542
rect -147 954 -89 966
rect -29 1542 29 1554
rect -29 966 -17 1542
rect 17 966 29 1542
rect -29 954 29 966
rect 89 1542 147 1554
rect 89 966 101 1542
rect 135 966 147 1542
rect 89 954 147 966
rect 207 1542 265 1554
rect 207 966 219 1542
rect 253 966 265 1542
rect 207 954 265 966
rect 325 1542 383 1554
rect 325 966 337 1542
rect 371 966 383 1542
rect 325 954 383 966
rect 443 1542 501 1554
rect 443 966 455 1542
rect 489 966 501 1542
rect 443 954 501 966
rect 561 1542 619 1554
rect 561 966 573 1542
rect 607 966 619 1542
rect 561 954 619 966
rect 679 1542 737 1554
rect 679 966 691 1542
rect 725 966 737 1542
rect 679 954 737 966
rect 797 1542 855 1554
rect 797 966 809 1542
rect 843 966 855 1542
rect 797 954 855 966
rect 915 1542 973 1554
rect 915 966 927 1542
rect 961 966 973 1542
rect 915 954 973 966
rect 1033 1542 1091 1554
rect 1033 966 1045 1542
rect 1079 966 1091 1542
rect 1033 954 1091 966
rect 1151 1542 1209 1554
rect 1151 966 1163 1542
rect 1197 966 1209 1542
rect 1151 954 1209 966
rect 1269 1542 1327 1554
rect 1269 966 1281 1542
rect 1315 966 1327 1542
rect 1269 954 1327 966
rect 1387 1542 1445 1554
rect 1387 966 1399 1542
rect 1433 966 1445 1542
rect 1387 954 1445 966
rect 1505 1542 1563 1554
rect 1505 966 1517 1542
rect 1551 966 1563 1542
rect 1505 954 1563 966
rect 1623 1542 1681 1554
rect 1623 966 1635 1542
rect 1669 966 1681 1542
rect 1623 954 1681 966
rect 1741 1542 1799 1554
rect 1741 966 1753 1542
rect 1787 966 1799 1542
rect 1741 954 1799 966
rect 1859 1542 1917 1554
rect 1859 966 1871 1542
rect 1905 966 1917 1542
rect 1859 954 1917 966
rect 1977 1542 2035 1554
rect 1977 966 1989 1542
rect 2023 966 2035 1542
rect 1977 954 2035 966
rect 2095 1542 2153 1554
rect 2095 966 2107 1542
rect 2141 966 2153 1542
rect 2095 954 2153 966
rect 2213 1542 2271 1554
rect 2213 966 2225 1542
rect 2259 966 2271 1542
rect 2213 954 2271 966
rect 2331 1542 2389 1554
rect 2331 966 2343 1542
rect 2377 966 2389 1542
rect 2331 954 2389 966
rect 2449 1542 2507 1554
rect 2449 966 2461 1542
rect 2495 966 2507 1542
rect 2449 954 2507 966
rect 2567 1542 2625 1554
rect 2567 966 2579 1542
rect 2613 966 2625 1542
rect 2567 954 2625 966
rect 2685 1542 2743 1554
rect 2685 966 2697 1542
rect 2731 966 2743 1542
rect 2685 954 2743 966
rect 2803 1542 2861 1554
rect 2803 966 2815 1542
rect 2849 966 2861 1542
rect 2803 954 2861 966
rect 2921 1542 2979 1554
rect 2921 966 2933 1542
rect 2967 966 2979 1542
rect 2921 954 2979 966
rect -2979 706 -2921 718
rect -2979 130 -2967 706
rect -2933 130 -2921 706
rect -2979 118 -2921 130
rect -2861 706 -2803 718
rect -2861 130 -2849 706
rect -2815 130 -2803 706
rect -2861 118 -2803 130
rect -2743 706 -2685 718
rect -2743 130 -2731 706
rect -2697 130 -2685 706
rect -2743 118 -2685 130
rect -2625 706 -2567 718
rect -2625 130 -2613 706
rect -2579 130 -2567 706
rect -2625 118 -2567 130
rect -2507 706 -2449 718
rect -2507 130 -2495 706
rect -2461 130 -2449 706
rect -2507 118 -2449 130
rect -2389 706 -2331 718
rect -2389 130 -2377 706
rect -2343 130 -2331 706
rect -2389 118 -2331 130
rect -2271 706 -2213 718
rect -2271 130 -2259 706
rect -2225 130 -2213 706
rect -2271 118 -2213 130
rect -2153 706 -2095 718
rect -2153 130 -2141 706
rect -2107 130 -2095 706
rect -2153 118 -2095 130
rect -2035 706 -1977 718
rect -2035 130 -2023 706
rect -1989 130 -1977 706
rect -2035 118 -1977 130
rect -1917 706 -1859 718
rect -1917 130 -1905 706
rect -1871 130 -1859 706
rect -1917 118 -1859 130
rect -1799 706 -1741 718
rect -1799 130 -1787 706
rect -1753 130 -1741 706
rect -1799 118 -1741 130
rect -1681 706 -1623 718
rect -1681 130 -1669 706
rect -1635 130 -1623 706
rect -1681 118 -1623 130
rect -1563 706 -1505 718
rect -1563 130 -1551 706
rect -1517 130 -1505 706
rect -1563 118 -1505 130
rect -1445 706 -1387 718
rect -1445 130 -1433 706
rect -1399 130 -1387 706
rect -1445 118 -1387 130
rect -1327 706 -1269 718
rect -1327 130 -1315 706
rect -1281 130 -1269 706
rect -1327 118 -1269 130
rect -1209 706 -1151 718
rect -1209 130 -1197 706
rect -1163 130 -1151 706
rect -1209 118 -1151 130
rect -1091 706 -1033 718
rect -1091 130 -1079 706
rect -1045 130 -1033 706
rect -1091 118 -1033 130
rect -973 706 -915 718
rect -973 130 -961 706
rect -927 130 -915 706
rect -973 118 -915 130
rect -855 706 -797 718
rect -855 130 -843 706
rect -809 130 -797 706
rect -855 118 -797 130
rect -737 706 -679 718
rect -737 130 -725 706
rect -691 130 -679 706
rect -737 118 -679 130
rect -619 706 -561 718
rect -619 130 -607 706
rect -573 130 -561 706
rect -619 118 -561 130
rect -501 706 -443 718
rect -501 130 -489 706
rect -455 130 -443 706
rect -501 118 -443 130
rect -383 706 -325 718
rect -383 130 -371 706
rect -337 130 -325 706
rect -383 118 -325 130
rect -265 706 -207 718
rect -265 130 -253 706
rect -219 130 -207 706
rect -265 118 -207 130
rect -147 706 -89 718
rect -147 130 -135 706
rect -101 130 -89 706
rect -147 118 -89 130
rect -29 706 29 718
rect -29 130 -17 706
rect 17 130 29 706
rect -29 118 29 130
rect 89 706 147 718
rect 89 130 101 706
rect 135 130 147 706
rect 89 118 147 130
rect 207 706 265 718
rect 207 130 219 706
rect 253 130 265 706
rect 207 118 265 130
rect 325 706 383 718
rect 325 130 337 706
rect 371 130 383 706
rect 325 118 383 130
rect 443 706 501 718
rect 443 130 455 706
rect 489 130 501 706
rect 443 118 501 130
rect 561 706 619 718
rect 561 130 573 706
rect 607 130 619 706
rect 561 118 619 130
rect 679 706 737 718
rect 679 130 691 706
rect 725 130 737 706
rect 679 118 737 130
rect 797 706 855 718
rect 797 130 809 706
rect 843 130 855 706
rect 797 118 855 130
rect 915 706 973 718
rect 915 130 927 706
rect 961 130 973 706
rect 915 118 973 130
rect 1033 706 1091 718
rect 1033 130 1045 706
rect 1079 130 1091 706
rect 1033 118 1091 130
rect 1151 706 1209 718
rect 1151 130 1163 706
rect 1197 130 1209 706
rect 1151 118 1209 130
rect 1269 706 1327 718
rect 1269 130 1281 706
rect 1315 130 1327 706
rect 1269 118 1327 130
rect 1387 706 1445 718
rect 1387 130 1399 706
rect 1433 130 1445 706
rect 1387 118 1445 130
rect 1505 706 1563 718
rect 1505 130 1517 706
rect 1551 130 1563 706
rect 1505 118 1563 130
rect 1623 706 1681 718
rect 1623 130 1635 706
rect 1669 130 1681 706
rect 1623 118 1681 130
rect 1741 706 1799 718
rect 1741 130 1753 706
rect 1787 130 1799 706
rect 1741 118 1799 130
rect 1859 706 1917 718
rect 1859 130 1871 706
rect 1905 130 1917 706
rect 1859 118 1917 130
rect 1977 706 2035 718
rect 1977 130 1989 706
rect 2023 130 2035 706
rect 1977 118 2035 130
rect 2095 706 2153 718
rect 2095 130 2107 706
rect 2141 130 2153 706
rect 2095 118 2153 130
rect 2213 706 2271 718
rect 2213 130 2225 706
rect 2259 130 2271 706
rect 2213 118 2271 130
rect 2331 706 2389 718
rect 2331 130 2343 706
rect 2377 130 2389 706
rect 2331 118 2389 130
rect 2449 706 2507 718
rect 2449 130 2461 706
rect 2495 130 2507 706
rect 2449 118 2507 130
rect 2567 706 2625 718
rect 2567 130 2579 706
rect 2613 130 2625 706
rect 2567 118 2625 130
rect 2685 706 2743 718
rect 2685 130 2697 706
rect 2731 130 2743 706
rect 2685 118 2743 130
rect 2803 706 2861 718
rect 2803 130 2815 706
rect 2849 130 2861 706
rect 2803 118 2861 130
rect 2921 706 2979 718
rect 2921 130 2933 706
rect 2967 130 2979 706
rect 2921 118 2979 130
rect -2979 -130 -2921 -118
rect -2979 -706 -2967 -130
rect -2933 -706 -2921 -130
rect -2979 -718 -2921 -706
rect -2861 -130 -2803 -118
rect -2861 -706 -2849 -130
rect -2815 -706 -2803 -130
rect -2861 -718 -2803 -706
rect -2743 -130 -2685 -118
rect -2743 -706 -2731 -130
rect -2697 -706 -2685 -130
rect -2743 -718 -2685 -706
rect -2625 -130 -2567 -118
rect -2625 -706 -2613 -130
rect -2579 -706 -2567 -130
rect -2625 -718 -2567 -706
rect -2507 -130 -2449 -118
rect -2507 -706 -2495 -130
rect -2461 -706 -2449 -130
rect -2507 -718 -2449 -706
rect -2389 -130 -2331 -118
rect -2389 -706 -2377 -130
rect -2343 -706 -2331 -130
rect -2389 -718 -2331 -706
rect -2271 -130 -2213 -118
rect -2271 -706 -2259 -130
rect -2225 -706 -2213 -130
rect -2271 -718 -2213 -706
rect -2153 -130 -2095 -118
rect -2153 -706 -2141 -130
rect -2107 -706 -2095 -130
rect -2153 -718 -2095 -706
rect -2035 -130 -1977 -118
rect -2035 -706 -2023 -130
rect -1989 -706 -1977 -130
rect -2035 -718 -1977 -706
rect -1917 -130 -1859 -118
rect -1917 -706 -1905 -130
rect -1871 -706 -1859 -130
rect -1917 -718 -1859 -706
rect -1799 -130 -1741 -118
rect -1799 -706 -1787 -130
rect -1753 -706 -1741 -130
rect -1799 -718 -1741 -706
rect -1681 -130 -1623 -118
rect -1681 -706 -1669 -130
rect -1635 -706 -1623 -130
rect -1681 -718 -1623 -706
rect -1563 -130 -1505 -118
rect -1563 -706 -1551 -130
rect -1517 -706 -1505 -130
rect -1563 -718 -1505 -706
rect -1445 -130 -1387 -118
rect -1445 -706 -1433 -130
rect -1399 -706 -1387 -130
rect -1445 -718 -1387 -706
rect -1327 -130 -1269 -118
rect -1327 -706 -1315 -130
rect -1281 -706 -1269 -130
rect -1327 -718 -1269 -706
rect -1209 -130 -1151 -118
rect -1209 -706 -1197 -130
rect -1163 -706 -1151 -130
rect -1209 -718 -1151 -706
rect -1091 -130 -1033 -118
rect -1091 -706 -1079 -130
rect -1045 -706 -1033 -130
rect -1091 -718 -1033 -706
rect -973 -130 -915 -118
rect -973 -706 -961 -130
rect -927 -706 -915 -130
rect -973 -718 -915 -706
rect -855 -130 -797 -118
rect -855 -706 -843 -130
rect -809 -706 -797 -130
rect -855 -718 -797 -706
rect -737 -130 -679 -118
rect -737 -706 -725 -130
rect -691 -706 -679 -130
rect -737 -718 -679 -706
rect -619 -130 -561 -118
rect -619 -706 -607 -130
rect -573 -706 -561 -130
rect -619 -718 -561 -706
rect -501 -130 -443 -118
rect -501 -706 -489 -130
rect -455 -706 -443 -130
rect -501 -718 -443 -706
rect -383 -130 -325 -118
rect -383 -706 -371 -130
rect -337 -706 -325 -130
rect -383 -718 -325 -706
rect -265 -130 -207 -118
rect -265 -706 -253 -130
rect -219 -706 -207 -130
rect -265 -718 -207 -706
rect -147 -130 -89 -118
rect -147 -706 -135 -130
rect -101 -706 -89 -130
rect -147 -718 -89 -706
rect -29 -130 29 -118
rect -29 -706 -17 -130
rect 17 -706 29 -130
rect -29 -718 29 -706
rect 89 -130 147 -118
rect 89 -706 101 -130
rect 135 -706 147 -130
rect 89 -718 147 -706
rect 207 -130 265 -118
rect 207 -706 219 -130
rect 253 -706 265 -130
rect 207 -718 265 -706
rect 325 -130 383 -118
rect 325 -706 337 -130
rect 371 -706 383 -130
rect 325 -718 383 -706
rect 443 -130 501 -118
rect 443 -706 455 -130
rect 489 -706 501 -130
rect 443 -718 501 -706
rect 561 -130 619 -118
rect 561 -706 573 -130
rect 607 -706 619 -130
rect 561 -718 619 -706
rect 679 -130 737 -118
rect 679 -706 691 -130
rect 725 -706 737 -130
rect 679 -718 737 -706
rect 797 -130 855 -118
rect 797 -706 809 -130
rect 843 -706 855 -130
rect 797 -718 855 -706
rect 915 -130 973 -118
rect 915 -706 927 -130
rect 961 -706 973 -130
rect 915 -718 973 -706
rect 1033 -130 1091 -118
rect 1033 -706 1045 -130
rect 1079 -706 1091 -130
rect 1033 -718 1091 -706
rect 1151 -130 1209 -118
rect 1151 -706 1163 -130
rect 1197 -706 1209 -130
rect 1151 -718 1209 -706
rect 1269 -130 1327 -118
rect 1269 -706 1281 -130
rect 1315 -706 1327 -130
rect 1269 -718 1327 -706
rect 1387 -130 1445 -118
rect 1387 -706 1399 -130
rect 1433 -706 1445 -130
rect 1387 -718 1445 -706
rect 1505 -130 1563 -118
rect 1505 -706 1517 -130
rect 1551 -706 1563 -130
rect 1505 -718 1563 -706
rect 1623 -130 1681 -118
rect 1623 -706 1635 -130
rect 1669 -706 1681 -130
rect 1623 -718 1681 -706
rect 1741 -130 1799 -118
rect 1741 -706 1753 -130
rect 1787 -706 1799 -130
rect 1741 -718 1799 -706
rect 1859 -130 1917 -118
rect 1859 -706 1871 -130
rect 1905 -706 1917 -130
rect 1859 -718 1917 -706
rect 1977 -130 2035 -118
rect 1977 -706 1989 -130
rect 2023 -706 2035 -130
rect 1977 -718 2035 -706
rect 2095 -130 2153 -118
rect 2095 -706 2107 -130
rect 2141 -706 2153 -130
rect 2095 -718 2153 -706
rect 2213 -130 2271 -118
rect 2213 -706 2225 -130
rect 2259 -706 2271 -130
rect 2213 -718 2271 -706
rect 2331 -130 2389 -118
rect 2331 -706 2343 -130
rect 2377 -706 2389 -130
rect 2331 -718 2389 -706
rect 2449 -130 2507 -118
rect 2449 -706 2461 -130
rect 2495 -706 2507 -130
rect 2449 -718 2507 -706
rect 2567 -130 2625 -118
rect 2567 -706 2579 -130
rect 2613 -706 2625 -130
rect 2567 -718 2625 -706
rect 2685 -130 2743 -118
rect 2685 -706 2697 -130
rect 2731 -706 2743 -130
rect 2685 -718 2743 -706
rect 2803 -130 2861 -118
rect 2803 -706 2815 -130
rect 2849 -706 2861 -130
rect 2803 -718 2861 -706
rect 2921 -130 2979 -118
rect 2921 -706 2933 -130
rect 2967 -706 2979 -130
rect 2921 -718 2979 -706
rect -2979 -966 -2921 -954
rect -2979 -1542 -2967 -966
rect -2933 -1542 -2921 -966
rect -2979 -1554 -2921 -1542
rect -2861 -966 -2803 -954
rect -2861 -1542 -2849 -966
rect -2815 -1542 -2803 -966
rect -2861 -1554 -2803 -1542
rect -2743 -966 -2685 -954
rect -2743 -1542 -2731 -966
rect -2697 -1542 -2685 -966
rect -2743 -1554 -2685 -1542
rect -2625 -966 -2567 -954
rect -2625 -1542 -2613 -966
rect -2579 -1542 -2567 -966
rect -2625 -1554 -2567 -1542
rect -2507 -966 -2449 -954
rect -2507 -1542 -2495 -966
rect -2461 -1542 -2449 -966
rect -2507 -1554 -2449 -1542
rect -2389 -966 -2331 -954
rect -2389 -1542 -2377 -966
rect -2343 -1542 -2331 -966
rect -2389 -1554 -2331 -1542
rect -2271 -966 -2213 -954
rect -2271 -1542 -2259 -966
rect -2225 -1542 -2213 -966
rect -2271 -1554 -2213 -1542
rect -2153 -966 -2095 -954
rect -2153 -1542 -2141 -966
rect -2107 -1542 -2095 -966
rect -2153 -1554 -2095 -1542
rect -2035 -966 -1977 -954
rect -2035 -1542 -2023 -966
rect -1989 -1542 -1977 -966
rect -2035 -1554 -1977 -1542
rect -1917 -966 -1859 -954
rect -1917 -1542 -1905 -966
rect -1871 -1542 -1859 -966
rect -1917 -1554 -1859 -1542
rect -1799 -966 -1741 -954
rect -1799 -1542 -1787 -966
rect -1753 -1542 -1741 -966
rect -1799 -1554 -1741 -1542
rect -1681 -966 -1623 -954
rect -1681 -1542 -1669 -966
rect -1635 -1542 -1623 -966
rect -1681 -1554 -1623 -1542
rect -1563 -966 -1505 -954
rect -1563 -1542 -1551 -966
rect -1517 -1542 -1505 -966
rect -1563 -1554 -1505 -1542
rect -1445 -966 -1387 -954
rect -1445 -1542 -1433 -966
rect -1399 -1542 -1387 -966
rect -1445 -1554 -1387 -1542
rect -1327 -966 -1269 -954
rect -1327 -1542 -1315 -966
rect -1281 -1542 -1269 -966
rect -1327 -1554 -1269 -1542
rect -1209 -966 -1151 -954
rect -1209 -1542 -1197 -966
rect -1163 -1542 -1151 -966
rect -1209 -1554 -1151 -1542
rect -1091 -966 -1033 -954
rect -1091 -1542 -1079 -966
rect -1045 -1542 -1033 -966
rect -1091 -1554 -1033 -1542
rect -973 -966 -915 -954
rect -973 -1542 -961 -966
rect -927 -1542 -915 -966
rect -973 -1554 -915 -1542
rect -855 -966 -797 -954
rect -855 -1542 -843 -966
rect -809 -1542 -797 -966
rect -855 -1554 -797 -1542
rect -737 -966 -679 -954
rect -737 -1542 -725 -966
rect -691 -1542 -679 -966
rect -737 -1554 -679 -1542
rect -619 -966 -561 -954
rect -619 -1542 -607 -966
rect -573 -1542 -561 -966
rect -619 -1554 -561 -1542
rect -501 -966 -443 -954
rect -501 -1542 -489 -966
rect -455 -1542 -443 -966
rect -501 -1554 -443 -1542
rect -383 -966 -325 -954
rect -383 -1542 -371 -966
rect -337 -1542 -325 -966
rect -383 -1554 -325 -1542
rect -265 -966 -207 -954
rect -265 -1542 -253 -966
rect -219 -1542 -207 -966
rect -265 -1554 -207 -1542
rect -147 -966 -89 -954
rect -147 -1542 -135 -966
rect -101 -1542 -89 -966
rect -147 -1554 -89 -1542
rect -29 -966 29 -954
rect -29 -1542 -17 -966
rect 17 -1542 29 -966
rect -29 -1554 29 -1542
rect 89 -966 147 -954
rect 89 -1542 101 -966
rect 135 -1542 147 -966
rect 89 -1554 147 -1542
rect 207 -966 265 -954
rect 207 -1542 219 -966
rect 253 -1542 265 -966
rect 207 -1554 265 -1542
rect 325 -966 383 -954
rect 325 -1542 337 -966
rect 371 -1542 383 -966
rect 325 -1554 383 -1542
rect 443 -966 501 -954
rect 443 -1542 455 -966
rect 489 -1542 501 -966
rect 443 -1554 501 -1542
rect 561 -966 619 -954
rect 561 -1542 573 -966
rect 607 -1542 619 -966
rect 561 -1554 619 -1542
rect 679 -966 737 -954
rect 679 -1542 691 -966
rect 725 -1542 737 -966
rect 679 -1554 737 -1542
rect 797 -966 855 -954
rect 797 -1542 809 -966
rect 843 -1542 855 -966
rect 797 -1554 855 -1542
rect 915 -966 973 -954
rect 915 -1542 927 -966
rect 961 -1542 973 -966
rect 915 -1554 973 -1542
rect 1033 -966 1091 -954
rect 1033 -1542 1045 -966
rect 1079 -1542 1091 -966
rect 1033 -1554 1091 -1542
rect 1151 -966 1209 -954
rect 1151 -1542 1163 -966
rect 1197 -1542 1209 -966
rect 1151 -1554 1209 -1542
rect 1269 -966 1327 -954
rect 1269 -1542 1281 -966
rect 1315 -1542 1327 -966
rect 1269 -1554 1327 -1542
rect 1387 -966 1445 -954
rect 1387 -1542 1399 -966
rect 1433 -1542 1445 -966
rect 1387 -1554 1445 -1542
rect 1505 -966 1563 -954
rect 1505 -1542 1517 -966
rect 1551 -1542 1563 -966
rect 1505 -1554 1563 -1542
rect 1623 -966 1681 -954
rect 1623 -1542 1635 -966
rect 1669 -1542 1681 -966
rect 1623 -1554 1681 -1542
rect 1741 -966 1799 -954
rect 1741 -1542 1753 -966
rect 1787 -1542 1799 -966
rect 1741 -1554 1799 -1542
rect 1859 -966 1917 -954
rect 1859 -1542 1871 -966
rect 1905 -1542 1917 -966
rect 1859 -1554 1917 -1542
rect 1977 -966 2035 -954
rect 1977 -1542 1989 -966
rect 2023 -1542 2035 -966
rect 1977 -1554 2035 -1542
rect 2095 -966 2153 -954
rect 2095 -1542 2107 -966
rect 2141 -1542 2153 -966
rect 2095 -1554 2153 -1542
rect 2213 -966 2271 -954
rect 2213 -1542 2225 -966
rect 2259 -1542 2271 -966
rect 2213 -1554 2271 -1542
rect 2331 -966 2389 -954
rect 2331 -1542 2343 -966
rect 2377 -1542 2389 -966
rect 2331 -1554 2389 -1542
rect 2449 -966 2507 -954
rect 2449 -1542 2461 -966
rect 2495 -1542 2507 -966
rect 2449 -1554 2507 -1542
rect 2567 -966 2625 -954
rect 2567 -1542 2579 -966
rect 2613 -1542 2625 -966
rect 2567 -1554 2625 -1542
rect 2685 -966 2743 -954
rect 2685 -1542 2697 -966
rect 2731 -1542 2743 -966
rect 2685 -1554 2743 -1542
rect 2803 -966 2861 -954
rect 2803 -1542 2815 -966
rect 2849 -1542 2861 -966
rect 2803 -1554 2861 -1542
rect 2921 -966 2979 -954
rect 2921 -1542 2933 -966
rect 2967 -1542 2979 -966
rect 2921 -1554 2979 -1542
<< pdiffc >>
rect -2967 966 -2933 1542
rect -2849 966 -2815 1542
rect -2731 966 -2697 1542
rect -2613 966 -2579 1542
rect -2495 966 -2461 1542
rect -2377 966 -2343 1542
rect -2259 966 -2225 1542
rect -2141 966 -2107 1542
rect -2023 966 -1989 1542
rect -1905 966 -1871 1542
rect -1787 966 -1753 1542
rect -1669 966 -1635 1542
rect -1551 966 -1517 1542
rect -1433 966 -1399 1542
rect -1315 966 -1281 1542
rect -1197 966 -1163 1542
rect -1079 966 -1045 1542
rect -961 966 -927 1542
rect -843 966 -809 1542
rect -725 966 -691 1542
rect -607 966 -573 1542
rect -489 966 -455 1542
rect -371 966 -337 1542
rect -253 966 -219 1542
rect -135 966 -101 1542
rect -17 966 17 1542
rect 101 966 135 1542
rect 219 966 253 1542
rect 337 966 371 1542
rect 455 966 489 1542
rect 573 966 607 1542
rect 691 966 725 1542
rect 809 966 843 1542
rect 927 966 961 1542
rect 1045 966 1079 1542
rect 1163 966 1197 1542
rect 1281 966 1315 1542
rect 1399 966 1433 1542
rect 1517 966 1551 1542
rect 1635 966 1669 1542
rect 1753 966 1787 1542
rect 1871 966 1905 1542
rect 1989 966 2023 1542
rect 2107 966 2141 1542
rect 2225 966 2259 1542
rect 2343 966 2377 1542
rect 2461 966 2495 1542
rect 2579 966 2613 1542
rect 2697 966 2731 1542
rect 2815 966 2849 1542
rect 2933 966 2967 1542
rect -2967 130 -2933 706
rect -2849 130 -2815 706
rect -2731 130 -2697 706
rect -2613 130 -2579 706
rect -2495 130 -2461 706
rect -2377 130 -2343 706
rect -2259 130 -2225 706
rect -2141 130 -2107 706
rect -2023 130 -1989 706
rect -1905 130 -1871 706
rect -1787 130 -1753 706
rect -1669 130 -1635 706
rect -1551 130 -1517 706
rect -1433 130 -1399 706
rect -1315 130 -1281 706
rect -1197 130 -1163 706
rect -1079 130 -1045 706
rect -961 130 -927 706
rect -843 130 -809 706
rect -725 130 -691 706
rect -607 130 -573 706
rect -489 130 -455 706
rect -371 130 -337 706
rect -253 130 -219 706
rect -135 130 -101 706
rect -17 130 17 706
rect 101 130 135 706
rect 219 130 253 706
rect 337 130 371 706
rect 455 130 489 706
rect 573 130 607 706
rect 691 130 725 706
rect 809 130 843 706
rect 927 130 961 706
rect 1045 130 1079 706
rect 1163 130 1197 706
rect 1281 130 1315 706
rect 1399 130 1433 706
rect 1517 130 1551 706
rect 1635 130 1669 706
rect 1753 130 1787 706
rect 1871 130 1905 706
rect 1989 130 2023 706
rect 2107 130 2141 706
rect 2225 130 2259 706
rect 2343 130 2377 706
rect 2461 130 2495 706
rect 2579 130 2613 706
rect 2697 130 2731 706
rect 2815 130 2849 706
rect 2933 130 2967 706
rect -2967 -706 -2933 -130
rect -2849 -706 -2815 -130
rect -2731 -706 -2697 -130
rect -2613 -706 -2579 -130
rect -2495 -706 -2461 -130
rect -2377 -706 -2343 -130
rect -2259 -706 -2225 -130
rect -2141 -706 -2107 -130
rect -2023 -706 -1989 -130
rect -1905 -706 -1871 -130
rect -1787 -706 -1753 -130
rect -1669 -706 -1635 -130
rect -1551 -706 -1517 -130
rect -1433 -706 -1399 -130
rect -1315 -706 -1281 -130
rect -1197 -706 -1163 -130
rect -1079 -706 -1045 -130
rect -961 -706 -927 -130
rect -843 -706 -809 -130
rect -725 -706 -691 -130
rect -607 -706 -573 -130
rect -489 -706 -455 -130
rect -371 -706 -337 -130
rect -253 -706 -219 -130
rect -135 -706 -101 -130
rect -17 -706 17 -130
rect 101 -706 135 -130
rect 219 -706 253 -130
rect 337 -706 371 -130
rect 455 -706 489 -130
rect 573 -706 607 -130
rect 691 -706 725 -130
rect 809 -706 843 -130
rect 927 -706 961 -130
rect 1045 -706 1079 -130
rect 1163 -706 1197 -130
rect 1281 -706 1315 -130
rect 1399 -706 1433 -130
rect 1517 -706 1551 -130
rect 1635 -706 1669 -130
rect 1753 -706 1787 -130
rect 1871 -706 1905 -130
rect 1989 -706 2023 -130
rect 2107 -706 2141 -130
rect 2225 -706 2259 -130
rect 2343 -706 2377 -130
rect 2461 -706 2495 -130
rect 2579 -706 2613 -130
rect 2697 -706 2731 -130
rect 2815 -706 2849 -130
rect 2933 -706 2967 -130
rect -2967 -1542 -2933 -966
rect -2849 -1542 -2815 -966
rect -2731 -1542 -2697 -966
rect -2613 -1542 -2579 -966
rect -2495 -1542 -2461 -966
rect -2377 -1542 -2343 -966
rect -2259 -1542 -2225 -966
rect -2141 -1542 -2107 -966
rect -2023 -1542 -1989 -966
rect -1905 -1542 -1871 -966
rect -1787 -1542 -1753 -966
rect -1669 -1542 -1635 -966
rect -1551 -1542 -1517 -966
rect -1433 -1542 -1399 -966
rect -1315 -1542 -1281 -966
rect -1197 -1542 -1163 -966
rect -1079 -1542 -1045 -966
rect -961 -1542 -927 -966
rect -843 -1542 -809 -966
rect -725 -1542 -691 -966
rect -607 -1542 -573 -966
rect -489 -1542 -455 -966
rect -371 -1542 -337 -966
rect -253 -1542 -219 -966
rect -135 -1542 -101 -966
rect -17 -1542 17 -966
rect 101 -1542 135 -966
rect 219 -1542 253 -966
rect 337 -1542 371 -966
rect 455 -1542 489 -966
rect 573 -1542 607 -966
rect 691 -1542 725 -966
rect 809 -1542 843 -966
rect 927 -1542 961 -966
rect 1045 -1542 1079 -966
rect 1163 -1542 1197 -966
rect 1281 -1542 1315 -966
rect 1399 -1542 1433 -966
rect 1517 -1542 1551 -966
rect 1635 -1542 1669 -966
rect 1753 -1542 1787 -966
rect 1871 -1542 1905 -966
rect 1989 -1542 2023 -966
rect 2107 -1542 2141 -966
rect 2225 -1542 2259 -966
rect 2343 -1542 2377 -966
rect 2461 -1542 2495 -966
rect 2579 -1542 2613 -966
rect 2697 -1542 2731 -966
rect 2815 -1542 2849 -966
rect 2933 -1542 2967 -966
<< nsubdiff >>
rect -3081 1703 -2985 1737
rect 2985 1703 3081 1737
rect -3081 1641 -3047 1703
rect 3047 1641 3081 1703
rect -3081 -1703 -3047 -1641
rect 3047 -1703 3081 -1641
rect -3081 -1737 -2985 -1703
rect 2985 -1737 3081 -1703
<< nsubdiffcont >>
rect -2985 1703 2985 1737
rect -3081 -1641 -3047 1641
rect 3047 -1641 3081 1641
rect -2985 -1737 2985 -1703
<< poly >>
rect -2924 1635 -2858 1651
rect -2924 1601 -2908 1635
rect -2874 1601 -2858 1635
rect -2924 1585 -2858 1601
rect -2806 1635 -2740 1651
rect -2806 1601 -2790 1635
rect -2756 1601 -2740 1635
rect -2806 1585 -2740 1601
rect -2688 1635 -2622 1651
rect -2688 1601 -2672 1635
rect -2638 1601 -2622 1635
rect -2688 1585 -2622 1601
rect -2570 1635 -2504 1651
rect -2570 1601 -2554 1635
rect -2520 1601 -2504 1635
rect -2570 1585 -2504 1601
rect -2452 1635 -2386 1651
rect -2452 1601 -2436 1635
rect -2402 1601 -2386 1635
rect -2452 1585 -2386 1601
rect -2334 1635 -2268 1651
rect -2334 1601 -2318 1635
rect -2284 1601 -2268 1635
rect -2334 1585 -2268 1601
rect -2216 1635 -2150 1651
rect -2216 1601 -2200 1635
rect -2166 1601 -2150 1635
rect -2216 1585 -2150 1601
rect -2098 1635 -2032 1651
rect -2098 1601 -2082 1635
rect -2048 1601 -2032 1635
rect -2098 1585 -2032 1601
rect -1980 1635 -1914 1651
rect -1980 1601 -1964 1635
rect -1930 1601 -1914 1635
rect -1980 1585 -1914 1601
rect -1862 1635 -1796 1651
rect -1862 1601 -1846 1635
rect -1812 1601 -1796 1635
rect -1862 1585 -1796 1601
rect -1744 1635 -1678 1651
rect -1744 1601 -1728 1635
rect -1694 1601 -1678 1635
rect -1744 1585 -1678 1601
rect -1626 1635 -1560 1651
rect -1626 1601 -1610 1635
rect -1576 1601 -1560 1635
rect -1626 1585 -1560 1601
rect -1508 1635 -1442 1651
rect -1508 1601 -1492 1635
rect -1458 1601 -1442 1635
rect -1508 1585 -1442 1601
rect -1390 1635 -1324 1651
rect -1390 1601 -1374 1635
rect -1340 1601 -1324 1635
rect -1390 1585 -1324 1601
rect -1272 1635 -1206 1651
rect -1272 1601 -1256 1635
rect -1222 1601 -1206 1635
rect -1272 1585 -1206 1601
rect -1154 1635 -1088 1651
rect -1154 1601 -1138 1635
rect -1104 1601 -1088 1635
rect -1154 1585 -1088 1601
rect -1036 1635 -970 1651
rect -1036 1601 -1020 1635
rect -986 1601 -970 1635
rect -1036 1585 -970 1601
rect -918 1635 -852 1651
rect -918 1601 -902 1635
rect -868 1601 -852 1635
rect -918 1585 -852 1601
rect -800 1635 -734 1651
rect -800 1601 -784 1635
rect -750 1601 -734 1635
rect -800 1585 -734 1601
rect -682 1635 -616 1651
rect -682 1601 -666 1635
rect -632 1601 -616 1635
rect -682 1585 -616 1601
rect -564 1635 -498 1651
rect -564 1601 -548 1635
rect -514 1601 -498 1635
rect -564 1585 -498 1601
rect -446 1635 -380 1651
rect -446 1601 -430 1635
rect -396 1601 -380 1635
rect -446 1585 -380 1601
rect -328 1635 -262 1651
rect -328 1601 -312 1635
rect -278 1601 -262 1635
rect -328 1585 -262 1601
rect -210 1635 -144 1651
rect -210 1601 -194 1635
rect -160 1601 -144 1635
rect -210 1585 -144 1601
rect -92 1635 -26 1651
rect -92 1601 -76 1635
rect -42 1601 -26 1635
rect -92 1585 -26 1601
rect 26 1635 92 1651
rect 26 1601 42 1635
rect 76 1601 92 1635
rect 26 1585 92 1601
rect 144 1635 210 1651
rect 144 1601 160 1635
rect 194 1601 210 1635
rect 144 1585 210 1601
rect 262 1635 328 1651
rect 262 1601 278 1635
rect 312 1601 328 1635
rect 262 1585 328 1601
rect 380 1635 446 1651
rect 380 1601 396 1635
rect 430 1601 446 1635
rect 380 1585 446 1601
rect 498 1635 564 1651
rect 498 1601 514 1635
rect 548 1601 564 1635
rect 498 1585 564 1601
rect 616 1635 682 1651
rect 616 1601 632 1635
rect 666 1601 682 1635
rect 616 1585 682 1601
rect 734 1635 800 1651
rect 734 1601 750 1635
rect 784 1601 800 1635
rect 734 1585 800 1601
rect 852 1635 918 1651
rect 852 1601 868 1635
rect 902 1601 918 1635
rect 852 1585 918 1601
rect 970 1635 1036 1651
rect 970 1601 986 1635
rect 1020 1601 1036 1635
rect 970 1585 1036 1601
rect 1088 1635 1154 1651
rect 1088 1601 1104 1635
rect 1138 1601 1154 1635
rect 1088 1585 1154 1601
rect 1206 1635 1272 1651
rect 1206 1601 1222 1635
rect 1256 1601 1272 1635
rect 1206 1585 1272 1601
rect 1324 1635 1390 1651
rect 1324 1601 1340 1635
rect 1374 1601 1390 1635
rect 1324 1585 1390 1601
rect 1442 1635 1508 1651
rect 1442 1601 1458 1635
rect 1492 1601 1508 1635
rect 1442 1585 1508 1601
rect 1560 1635 1626 1651
rect 1560 1601 1576 1635
rect 1610 1601 1626 1635
rect 1560 1585 1626 1601
rect 1678 1635 1744 1651
rect 1678 1601 1694 1635
rect 1728 1601 1744 1635
rect 1678 1585 1744 1601
rect 1796 1635 1862 1651
rect 1796 1601 1812 1635
rect 1846 1601 1862 1635
rect 1796 1585 1862 1601
rect 1914 1635 1980 1651
rect 1914 1601 1930 1635
rect 1964 1601 1980 1635
rect 1914 1585 1980 1601
rect 2032 1635 2098 1651
rect 2032 1601 2048 1635
rect 2082 1601 2098 1635
rect 2032 1585 2098 1601
rect 2150 1635 2216 1651
rect 2150 1601 2166 1635
rect 2200 1601 2216 1635
rect 2150 1585 2216 1601
rect 2268 1635 2334 1651
rect 2268 1601 2284 1635
rect 2318 1601 2334 1635
rect 2268 1585 2334 1601
rect 2386 1635 2452 1651
rect 2386 1601 2402 1635
rect 2436 1601 2452 1635
rect 2386 1585 2452 1601
rect 2504 1635 2570 1651
rect 2504 1601 2520 1635
rect 2554 1601 2570 1635
rect 2504 1585 2570 1601
rect 2622 1635 2688 1651
rect 2622 1601 2638 1635
rect 2672 1601 2688 1635
rect 2622 1585 2688 1601
rect 2740 1635 2806 1651
rect 2740 1601 2756 1635
rect 2790 1601 2806 1635
rect 2740 1585 2806 1601
rect 2858 1635 2924 1651
rect 2858 1601 2874 1635
rect 2908 1601 2924 1635
rect 2858 1585 2924 1601
rect -2921 1554 -2861 1585
rect -2803 1554 -2743 1585
rect -2685 1554 -2625 1585
rect -2567 1554 -2507 1585
rect -2449 1554 -2389 1585
rect -2331 1554 -2271 1585
rect -2213 1554 -2153 1585
rect -2095 1554 -2035 1585
rect -1977 1554 -1917 1585
rect -1859 1554 -1799 1585
rect -1741 1554 -1681 1585
rect -1623 1554 -1563 1585
rect -1505 1554 -1445 1585
rect -1387 1554 -1327 1585
rect -1269 1554 -1209 1585
rect -1151 1554 -1091 1585
rect -1033 1554 -973 1585
rect -915 1554 -855 1585
rect -797 1554 -737 1585
rect -679 1554 -619 1585
rect -561 1554 -501 1585
rect -443 1554 -383 1585
rect -325 1554 -265 1585
rect -207 1554 -147 1585
rect -89 1554 -29 1585
rect 29 1554 89 1585
rect 147 1554 207 1585
rect 265 1554 325 1585
rect 383 1554 443 1585
rect 501 1554 561 1585
rect 619 1554 679 1585
rect 737 1554 797 1585
rect 855 1554 915 1585
rect 973 1554 1033 1585
rect 1091 1554 1151 1585
rect 1209 1554 1269 1585
rect 1327 1554 1387 1585
rect 1445 1554 1505 1585
rect 1563 1554 1623 1585
rect 1681 1554 1741 1585
rect 1799 1554 1859 1585
rect 1917 1554 1977 1585
rect 2035 1554 2095 1585
rect 2153 1554 2213 1585
rect 2271 1554 2331 1585
rect 2389 1554 2449 1585
rect 2507 1554 2567 1585
rect 2625 1554 2685 1585
rect 2743 1554 2803 1585
rect 2861 1554 2921 1585
rect -2921 923 -2861 954
rect -2803 923 -2743 954
rect -2685 923 -2625 954
rect -2567 923 -2507 954
rect -2449 923 -2389 954
rect -2331 923 -2271 954
rect -2213 923 -2153 954
rect -2095 923 -2035 954
rect -1977 923 -1917 954
rect -1859 923 -1799 954
rect -1741 923 -1681 954
rect -1623 923 -1563 954
rect -1505 923 -1445 954
rect -1387 923 -1327 954
rect -1269 923 -1209 954
rect -1151 923 -1091 954
rect -1033 923 -973 954
rect -915 923 -855 954
rect -797 923 -737 954
rect -679 923 -619 954
rect -561 923 -501 954
rect -443 923 -383 954
rect -325 923 -265 954
rect -207 923 -147 954
rect -89 923 -29 954
rect 29 923 89 954
rect 147 923 207 954
rect 265 923 325 954
rect 383 923 443 954
rect 501 923 561 954
rect 619 923 679 954
rect 737 923 797 954
rect 855 923 915 954
rect 973 923 1033 954
rect 1091 923 1151 954
rect 1209 923 1269 954
rect 1327 923 1387 954
rect 1445 923 1505 954
rect 1563 923 1623 954
rect 1681 923 1741 954
rect 1799 923 1859 954
rect 1917 923 1977 954
rect 2035 923 2095 954
rect 2153 923 2213 954
rect 2271 923 2331 954
rect 2389 923 2449 954
rect 2507 923 2567 954
rect 2625 923 2685 954
rect 2743 923 2803 954
rect 2861 923 2921 954
rect -2924 907 -2858 923
rect -2924 873 -2908 907
rect -2874 873 -2858 907
rect -2924 857 -2858 873
rect -2806 907 -2740 923
rect -2806 873 -2790 907
rect -2756 873 -2740 907
rect -2806 857 -2740 873
rect -2688 907 -2622 923
rect -2688 873 -2672 907
rect -2638 873 -2622 907
rect -2688 857 -2622 873
rect -2570 907 -2504 923
rect -2570 873 -2554 907
rect -2520 873 -2504 907
rect -2570 857 -2504 873
rect -2452 907 -2386 923
rect -2452 873 -2436 907
rect -2402 873 -2386 907
rect -2452 857 -2386 873
rect -2334 907 -2268 923
rect -2334 873 -2318 907
rect -2284 873 -2268 907
rect -2334 857 -2268 873
rect -2216 907 -2150 923
rect -2216 873 -2200 907
rect -2166 873 -2150 907
rect -2216 857 -2150 873
rect -2098 907 -2032 923
rect -2098 873 -2082 907
rect -2048 873 -2032 907
rect -2098 857 -2032 873
rect -1980 907 -1914 923
rect -1980 873 -1964 907
rect -1930 873 -1914 907
rect -1980 857 -1914 873
rect -1862 907 -1796 923
rect -1862 873 -1846 907
rect -1812 873 -1796 907
rect -1862 857 -1796 873
rect -1744 907 -1678 923
rect -1744 873 -1728 907
rect -1694 873 -1678 907
rect -1744 857 -1678 873
rect -1626 907 -1560 923
rect -1626 873 -1610 907
rect -1576 873 -1560 907
rect -1626 857 -1560 873
rect -1508 907 -1442 923
rect -1508 873 -1492 907
rect -1458 873 -1442 907
rect -1508 857 -1442 873
rect -1390 907 -1324 923
rect -1390 873 -1374 907
rect -1340 873 -1324 907
rect -1390 857 -1324 873
rect -1272 907 -1206 923
rect -1272 873 -1256 907
rect -1222 873 -1206 907
rect -1272 857 -1206 873
rect -1154 907 -1088 923
rect -1154 873 -1138 907
rect -1104 873 -1088 907
rect -1154 857 -1088 873
rect -1036 907 -970 923
rect -1036 873 -1020 907
rect -986 873 -970 907
rect -1036 857 -970 873
rect -918 907 -852 923
rect -918 873 -902 907
rect -868 873 -852 907
rect -918 857 -852 873
rect -800 907 -734 923
rect -800 873 -784 907
rect -750 873 -734 907
rect -800 857 -734 873
rect -682 907 -616 923
rect -682 873 -666 907
rect -632 873 -616 907
rect -682 857 -616 873
rect -564 907 -498 923
rect -564 873 -548 907
rect -514 873 -498 907
rect -564 857 -498 873
rect -446 907 -380 923
rect -446 873 -430 907
rect -396 873 -380 907
rect -446 857 -380 873
rect -328 907 -262 923
rect -328 873 -312 907
rect -278 873 -262 907
rect -328 857 -262 873
rect -210 907 -144 923
rect -210 873 -194 907
rect -160 873 -144 907
rect -210 857 -144 873
rect -92 907 -26 923
rect -92 873 -76 907
rect -42 873 -26 907
rect -92 857 -26 873
rect 26 907 92 923
rect 26 873 42 907
rect 76 873 92 907
rect 26 857 92 873
rect 144 907 210 923
rect 144 873 160 907
rect 194 873 210 907
rect 144 857 210 873
rect 262 907 328 923
rect 262 873 278 907
rect 312 873 328 907
rect 262 857 328 873
rect 380 907 446 923
rect 380 873 396 907
rect 430 873 446 907
rect 380 857 446 873
rect 498 907 564 923
rect 498 873 514 907
rect 548 873 564 907
rect 498 857 564 873
rect 616 907 682 923
rect 616 873 632 907
rect 666 873 682 907
rect 616 857 682 873
rect 734 907 800 923
rect 734 873 750 907
rect 784 873 800 907
rect 734 857 800 873
rect 852 907 918 923
rect 852 873 868 907
rect 902 873 918 907
rect 852 857 918 873
rect 970 907 1036 923
rect 970 873 986 907
rect 1020 873 1036 907
rect 970 857 1036 873
rect 1088 907 1154 923
rect 1088 873 1104 907
rect 1138 873 1154 907
rect 1088 857 1154 873
rect 1206 907 1272 923
rect 1206 873 1222 907
rect 1256 873 1272 907
rect 1206 857 1272 873
rect 1324 907 1390 923
rect 1324 873 1340 907
rect 1374 873 1390 907
rect 1324 857 1390 873
rect 1442 907 1508 923
rect 1442 873 1458 907
rect 1492 873 1508 907
rect 1442 857 1508 873
rect 1560 907 1626 923
rect 1560 873 1576 907
rect 1610 873 1626 907
rect 1560 857 1626 873
rect 1678 907 1744 923
rect 1678 873 1694 907
rect 1728 873 1744 907
rect 1678 857 1744 873
rect 1796 907 1862 923
rect 1796 873 1812 907
rect 1846 873 1862 907
rect 1796 857 1862 873
rect 1914 907 1980 923
rect 1914 873 1930 907
rect 1964 873 1980 907
rect 1914 857 1980 873
rect 2032 907 2098 923
rect 2032 873 2048 907
rect 2082 873 2098 907
rect 2032 857 2098 873
rect 2150 907 2216 923
rect 2150 873 2166 907
rect 2200 873 2216 907
rect 2150 857 2216 873
rect 2268 907 2334 923
rect 2268 873 2284 907
rect 2318 873 2334 907
rect 2268 857 2334 873
rect 2386 907 2452 923
rect 2386 873 2402 907
rect 2436 873 2452 907
rect 2386 857 2452 873
rect 2504 907 2570 923
rect 2504 873 2520 907
rect 2554 873 2570 907
rect 2504 857 2570 873
rect 2622 907 2688 923
rect 2622 873 2638 907
rect 2672 873 2688 907
rect 2622 857 2688 873
rect 2740 907 2806 923
rect 2740 873 2756 907
rect 2790 873 2806 907
rect 2740 857 2806 873
rect 2858 907 2924 923
rect 2858 873 2874 907
rect 2908 873 2924 907
rect 2858 857 2924 873
rect -2924 799 -2858 815
rect -2924 765 -2908 799
rect -2874 765 -2858 799
rect -2924 749 -2858 765
rect -2806 799 -2740 815
rect -2806 765 -2790 799
rect -2756 765 -2740 799
rect -2806 749 -2740 765
rect -2688 799 -2622 815
rect -2688 765 -2672 799
rect -2638 765 -2622 799
rect -2688 749 -2622 765
rect -2570 799 -2504 815
rect -2570 765 -2554 799
rect -2520 765 -2504 799
rect -2570 749 -2504 765
rect -2452 799 -2386 815
rect -2452 765 -2436 799
rect -2402 765 -2386 799
rect -2452 749 -2386 765
rect -2334 799 -2268 815
rect -2334 765 -2318 799
rect -2284 765 -2268 799
rect -2334 749 -2268 765
rect -2216 799 -2150 815
rect -2216 765 -2200 799
rect -2166 765 -2150 799
rect -2216 749 -2150 765
rect -2098 799 -2032 815
rect -2098 765 -2082 799
rect -2048 765 -2032 799
rect -2098 749 -2032 765
rect -1980 799 -1914 815
rect -1980 765 -1964 799
rect -1930 765 -1914 799
rect -1980 749 -1914 765
rect -1862 799 -1796 815
rect -1862 765 -1846 799
rect -1812 765 -1796 799
rect -1862 749 -1796 765
rect -1744 799 -1678 815
rect -1744 765 -1728 799
rect -1694 765 -1678 799
rect -1744 749 -1678 765
rect -1626 799 -1560 815
rect -1626 765 -1610 799
rect -1576 765 -1560 799
rect -1626 749 -1560 765
rect -1508 799 -1442 815
rect -1508 765 -1492 799
rect -1458 765 -1442 799
rect -1508 749 -1442 765
rect -1390 799 -1324 815
rect -1390 765 -1374 799
rect -1340 765 -1324 799
rect -1390 749 -1324 765
rect -1272 799 -1206 815
rect -1272 765 -1256 799
rect -1222 765 -1206 799
rect -1272 749 -1206 765
rect -1154 799 -1088 815
rect -1154 765 -1138 799
rect -1104 765 -1088 799
rect -1154 749 -1088 765
rect -1036 799 -970 815
rect -1036 765 -1020 799
rect -986 765 -970 799
rect -1036 749 -970 765
rect -918 799 -852 815
rect -918 765 -902 799
rect -868 765 -852 799
rect -918 749 -852 765
rect -800 799 -734 815
rect -800 765 -784 799
rect -750 765 -734 799
rect -800 749 -734 765
rect -682 799 -616 815
rect -682 765 -666 799
rect -632 765 -616 799
rect -682 749 -616 765
rect -564 799 -498 815
rect -564 765 -548 799
rect -514 765 -498 799
rect -564 749 -498 765
rect -446 799 -380 815
rect -446 765 -430 799
rect -396 765 -380 799
rect -446 749 -380 765
rect -328 799 -262 815
rect -328 765 -312 799
rect -278 765 -262 799
rect -328 749 -262 765
rect -210 799 -144 815
rect -210 765 -194 799
rect -160 765 -144 799
rect -210 749 -144 765
rect -92 799 -26 815
rect -92 765 -76 799
rect -42 765 -26 799
rect -92 749 -26 765
rect 26 799 92 815
rect 26 765 42 799
rect 76 765 92 799
rect 26 749 92 765
rect 144 799 210 815
rect 144 765 160 799
rect 194 765 210 799
rect 144 749 210 765
rect 262 799 328 815
rect 262 765 278 799
rect 312 765 328 799
rect 262 749 328 765
rect 380 799 446 815
rect 380 765 396 799
rect 430 765 446 799
rect 380 749 446 765
rect 498 799 564 815
rect 498 765 514 799
rect 548 765 564 799
rect 498 749 564 765
rect 616 799 682 815
rect 616 765 632 799
rect 666 765 682 799
rect 616 749 682 765
rect 734 799 800 815
rect 734 765 750 799
rect 784 765 800 799
rect 734 749 800 765
rect 852 799 918 815
rect 852 765 868 799
rect 902 765 918 799
rect 852 749 918 765
rect 970 799 1036 815
rect 970 765 986 799
rect 1020 765 1036 799
rect 970 749 1036 765
rect 1088 799 1154 815
rect 1088 765 1104 799
rect 1138 765 1154 799
rect 1088 749 1154 765
rect 1206 799 1272 815
rect 1206 765 1222 799
rect 1256 765 1272 799
rect 1206 749 1272 765
rect 1324 799 1390 815
rect 1324 765 1340 799
rect 1374 765 1390 799
rect 1324 749 1390 765
rect 1442 799 1508 815
rect 1442 765 1458 799
rect 1492 765 1508 799
rect 1442 749 1508 765
rect 1560 799 1626 815
rect 1560 765 1576 799
rect 1610 765 1626 799
rect 1560 749 1626 765
rect 1678 799 1744 815
rect 1678 765 1694 799
rect 1728 765 1744 799
rect 1678 749 1744 765
rect 1796 799 1862 815
rect 1796 765 1812 799
rect 1846 765 1862 799
rect 1796 749 1862 765
rect 1914 799 1980 815
rect 1914 765 1930 799
rect 1964 765 1980 799
rect 1914 749 1980 765
rect 2032 799 2098 815
rect 2032 765 2048 799
rect 2082 765 2098 799
rect 2032 749 2098 765
rect 2150 799 2216 815
rect 2150 765 2166 799
rect 2200 765 2216 799
rect 2150 749 2216 765
rect 2268 799 2334 815
rect 2268 765 2284 799
rect 2318 765 2334 799
rect 2268 749 2334 765
rect 2386 799 2452 815
rect 2386 765 2402 799
rect 2436 765 2452 799
rect 2386 749 2452 765
rect 2504 799 2570 815
rect 2504 765 2520 799
rect 2554 765 2570 799
rect 2504 749 2570 765
rect 2622 799 2688 815
rect 2622 765 2638 799
rect 2672 765 2688 799
rect 2622 749 2688 765
rect 2740 799 2806 815
rect 2740 765 2756 799
rect 2790 765 2806 799
rect 2740 749 2806 765
rect 2858 799 2924 815
rect 2858 765 2874 799
rect 2908 765 2924 799
rect 2858 749 2924 765
rect -2921 718 -2861 749
rect -2803 718 -2743 749
rect -2685 718 -2625 749
rect -2567 718 -2507 749
rect -2449 718 -2389 749
rect -2331 718 -2271 749
rect -2213 718 -2153 749
rect -2095 718 -2035 749
rect -1977 718 -1917 749
rect -1859 718 -1799 749
rect -1741 718 -1681 749
rect -1623 718 -1563 749
rect -1505 718 -1445 749
rect -1387 718 -1327 749
rect -1269 718 -1209 749
rect -1151 718 -1091 749
rect -1033 718 -973 749
rect -915 718 -855 749
rect -797 718 -737 749
rect -679 718 -619 749
rect -561 718 -501 749
rect -443 718 -383 749
rect -325 718 -265 749
rect -207 718 -147 749
rect -89 718 -29 749
rect 29 718 89 749
rect 147 718 207 749
rect 265 718 325 749
rect 383 718 443 749
rect 501 718 561 749
rect 619 718 679 749
rect 737 718 797 749
rect 855 718 915 749
rect 973 718 1033 749
rect 1091 718 1151 749
rect 1209 718 1269 749
rect 1327 718 1387 749
rect 1445 718 1505 749
rect 1563 718 1623 749
rect 1681 718 1741 749
rect 1799 718 1859 749
rect 1917 718 1977 749
rect 2035 718 2095 749
rect 2153 718 2213 749
rect 2271 718 2331 749
rect 2389 718 2449 749
rect 2507 718 2567 749
rect 2625 718 2685 749
rect 2743 718 2803 749
rect 2861 718 2921 749
rect -2921 87 -2861 118
rect -2803 87 -2743 118
rect -2685 87 -2625 118
rect -2567 87 -2507 118
rect -2449 87 -2389 118
rect -2331 87 -2271 118
rect -2213 87 -2153 118
rect -2095 87 -2035 118
rect -1977 87 -1917 118
rect -1859 87 -1799 118
rect -1741 87 -1681 118
rect -1623 87 -1563 118
rect -1505 87 -1445 118
rect -1387 87 -1327 118
rect -1269 87 -1209 118
rect -1151 87 -1091 118
rect -1033 87 -973 118
rect -915 87 -855 118
rect -797 87 -737 118
rect -679 87 -619 118
rect -561 87 -501 118
rect -443 87 -383 118
rect -325 87 -265 118
rect -207 87 -147 118
rect -89 87 -29 118
rect 29 87 89 118
rect 147 87 207 118
rect 265 87 325 118
rect 383 87 443 118
rect 501 87 561 118
rect 619 87 679 118
rect 737 87 797 118
rect 855 87 915 118
rect 973 87 1033 118
rect 1091 87 1151 118
rect 1209 87 1269 118
rect 1327 87 1387 118
rect 1445 87 1505 118
rect 1563 87 1623 118
rect 1681 87 1741 118
rect 1799 87 1859 118
rect 1917 87 1977 118
rect 2035 87 2095 118
rect 2153 87 2213 118
rect 2271 87 2331 118
rect 2389 87 2449 118
rect 2507 87 2567 118
rect 2625 87 2685 118
rect 2743 87 2803 118
rect 2861 87 2921 118
rect -2924 71 -2858 87
rect -2924 37 -2908 71
rect -2874 37 -2858 71
rect -2924 21 -2858 37
rect -2806 71 -2740 87
rect -2806 37 -2790 71
rect -2756 37 -2740 71
rect -2806 21 -2740 37
rect -2688 71 -2622 87
rect -2688 37 -2672 71
rect -2638 37 -2622 71
rect -2688 21 -2622 37
rect -2570 71 -2504 87
rect -2570 37 -2554 71
rect -2520 37 -2504 71
rect -2570 21 -2504 37
rect -2452 71 -2386 87
rect -2452 37 -2436 71
rect -2402 37 -2386 71
rect -2452 21 -2386 37
rect -2334 71 -2268 87
rect -2334 37 -2318 71
rect -2284 37 -2268 71
rect -2334 21 -2268 37
rect -2216 71 -2150 87
rect -2216 37 -2200 71
rect -2166 37 -2150 71
rect -2216 21 -2150 37
rect -2098 71 -2032 87
rect -2098 37 -2082 71
rect -2048 37 -2032 71
rect -2098 21 -2032 37
rect -1980 71 -1914 87
rect -1980 37 -1964 71
rect -1930 37 -1914 71
rect -1980 21 -1914 37
rect -1862 71 -1796 87
rect -1862 37 -1846 71
rect -1812 37 -1796 71
rect -1862 21 -1796 37
rect -1744 71 -1678 87
rect -1744 37 -1728 71
rect -1694 37 -1678 71
rect -1744 21 -1678 37
rect -1626 71 -1560 87
rect -1626 37 -1610 71
rect -1576 37 -1560 71
rect -1626 21 -1560 37
rect -1508 71 -1442 87
rect -1508 37 -1492 71
rect -1458 37 -1442 71
rect -1508 21 -1442 37
rect -1390 71 -1324 87
rect -1390 37 -1374 71
rect -1340 37 -1324 71
rect -1390 21 -1324 37
rect -1272 71 -1206 87
rect -1272 37 -1256 71
rect -1222 37 -1206 71
rect -1272 21 -1206 37
rect -1154 71 -1088 87
rect -1154 37 -1138 71
rect -1104 37 -1088 71
rect -1154 21 -1088 37
rect -1036 71 -970 87
rect -1036 37 -1020 71
rect -986 37 -970 71
rect -1036 21 -970 37
rect -918 71 -852 87
rect -918 37 -902 71
rect -868 37 -852 71
rect -918 21 -852 37
rect -800 71 -734 87
rect -800 37 -784 71
rect -750 37 -734 71
rect -800 21 -734 37
rect -682 71 -616 87
rect -682 37 -666 71
rect -632 37 -616 71
rect -682 21 -616 37
rect -564 71 -498 87
rect -564 37 -548 71
rect -514 37 -498 71
rect -564 21 -498 37
rect -446 71 -380 87
rect -446 37 -430 71
rect -396 37 -380 71
rect -446 21 -380 37
rect -328 71 -262 87
rect -328 37 -312 71
rect -278 37 -262 71
rect -328 21 -262 37
rect -210 71 -144 87
rect -210 37 -194 71
rect -160 37 -144 71
rect -210 21 -144 37
rect -92 71 -26 87
rect -92 37 -76 71
rect -42 37 -26 71
rect -92 21 -26 37
rect 26 71 92 87
rect 26 37 42 71
rect 76 37 92 71
rect 26 21 92 37
rect 144 71 210 87
rect 144 37 160 71
rect 194 37 210 71
rect 144 21 210 37
rect 262 71 328 87
rect 262 37 278 71
rect 312 37 328 71
rect 262 21 328 37
rect 380 71 446 87
rect 380 37 396 71
rect 430 37 446 71
rect 380 21 446 37
rect 498 71 564 87
rect 498 37 514 71
rect 548 37 564 71
rect 498 21 564 37
rect 616 71 682 87
rect 616 37 632 71
rect 666 37 682 71
rect 616 21 682 37
rect 734 71 800 87
rect 734 37 750 71
rect 784 37 800 71
rect 734 21 800 37
rect 852 71 918 87
rect 852 37 868 71
rect 902 37 918 71
rect 852 21 918 37
rect 970 71 1036 87
rect 970 37 986 71
rect 1020 37 1036 71
rect 970 21 1036 37
rect 1088 71 1154 87
rect 1088 37 1104 71
rect 1138 37 1154 71
rect 1088 21 1154 37
rect 1206 71 1272 87
rect 1206 37 1222 71
rect 1256 37 1272 71
rect 1206 21 1272 37
rect 1324 71 1390 87
rect 1324 37 1340 71
rect 1374 37 1390 71
rect 1324 21 1390 37
rect 1442 71 1508 87
rect 1442 37 1458 71
rect 1492 37 1508 71
rect 1442 21 1508 37
rect 1560 71 1626 87
rect 1560 37 1576 71
rect 1610 37 1626 71
rect 1560 21 1626 37
rect 1678 71 1744 87
rect 1678 37 1694 71
rect 1728 37 1744 71
rect 1678 21 1744 37
rect 1796 71 1862 87
rect 1796 37 1812 71
rect 1846 37 1862 71
rect 1796 21 1862 37
rect 1914 71 1980 87
rect 1914 37 1930 71
rect 1964 37 1980 71
rect 1914 21 1980 37
rect 2032 71 2098 87
rect 2032 37 2048 71
rect 2082 37 2098 71
rect 2032 21 2098 37
rect 2150 71 2216 87
rect 2150 37 2166 71
rect 2200 37 2216 71
rect 2150 21 2216 37
rect 2268 71 2334 87
rect 2268 37 2284 71
rect 2318 37 2334 71
rect 2268 21 2334 37
rect 2386 71 2452 87
rect 2386 37 2402 71
rect 2436 37 2452 71
rect 2386 21 2452 37
rect 2504 71 2570 87
rect 2504 37 2520 71
rect 2554 37 2570 71
rect 2504 21 2570 37
rect 2622 71 2688 87
rect 2622 37 2638 71
rect 2672 37 2688 71
rect 2622 21 2688 37
rect 2740 71 2806 87
rect 2740 37 2756 71
rect 2790 37 2806 71
rect 2740 21 2806 37
rect 2858 71 2924 87
rect 2858 37 2874 71
rect 2908 37 2924 71
rect 2858 21 2924 37
rect -2924 -37 -2858 -21
rect -2924 -71 -2908 -37
rect -2874 -71 -2858 -37
rect -2924 -87 -2858 -71
rect -2806 -37 -2740 -21
rect -2806 -71 -2790 -37
rect -2756 -71 -2740 -37
rect -2806 -87 -2740 -71
rect -2688 -37 -2622 -21
rect -2688 -71 -2672 -37
rect -2638 -71 -2622 -37
rect -2688 -87 -2622 -71
rect -2570 -37 -2504 -21
rect -2570 -71 -2554 -37
rect -2520 -71 -2504 -37
rect -2570 -87 -2504 -71
rect -2452 -37 -2386 -21
rect -2452 -71 -2436 -37
rect -2402 -71 -2386 -37
rect -2452 -87 -2386 -71
rect -2334 -37 -2268 -21
rect -2334 -71 -2318 -37
rect -2284 -71 -2268 -37
rect -2334 -87 -2268 -71
rect -2216 -37 -2150 -21
rect -2216 -71 -2200 -37
rect -2166 -71 -2150 -37
rect -2216 -87 -2150 -71
rect -2098 -37 -2032 -21
rect -2098 -71 -2082 -37
rect -2048 -71 -2032 -37
rect -2098 -87 -2032 -71
rect -1980 -37 -1914 -21
rect -1980 -71 -1964 -37
rect -1930 -71 -1914 -37
rect -1980 -87 -1914 -71
rect -1862 -37 -1796 -21
rect -1862 -71 -1846 -37
rect -1812 -71 -1796 -37
rect -1862 -87 -1796 -71
rect -1744 -37 -1678 -21
rect -1744 -71 -1728 -37
rect -1694 -71 -1678 -37
rect -1744 -87 -1678 -71
rect -1626 -37 -1560 -21
rect -1626 -71 -1610 -37
rect -1576 -71 -1560 -37
rect -1626 -87 -1560 -71
rect -1508 -37 -1442 -21
rect -1508 -71 -1492 -37
rect -1458 -71 -1442 -37
rect -1508 -87 -1442 -71
rect -1390 -37 -1324 -21
rect -1390 -71 -1374 -37
rect -1340 -71 -1324 -37
rect -1390 -87 -1324 -71
rect -1272 -37 -1206 -21
rect -1272 -71 -1256 -37
rect -1222 -71 -1206 -37
rect -1272 -87 -1206 -71
rect -1154 -37 -1088 -21
rect -1154 -71 -1138 -37
rect -1104 -71 -1088 -37
rect -1154 -87 -1088 -71
rect -1036 -37 -970 -21
rect -1036 -71 -1020 -37
rect -986 -71 -970 -37
rect -1036 -87 -970 -71
rect -918 -37 -852 -21
rect -918 -71 -902 -37
rect -868 -71 -852 -37
rect -918 -87 -852 -71
rect -800 -37 -734 -21
rect -800 -71 -784 -37
rect -750 -71 -734 -37
rect -800 -87 -734 -71
rect -682 -37 -616 -21
rect -682 -71 -666 -37
rect -632 -71 -616 -37
rect -682 -87 -616 -71
rect -564 -37 -498 -21
rect -564 -71 -548 -37
rect -514 -71 -498 -37
rect -564 -87 -498 -71
rect -446 -37 -380 -21
rect -446 -71 -430 -37
rect -396 -71 -380 -37
rect -446 -87 -380 -71
rect -328 -37 -262 -21
rect -328 -71 -312 -37
rect -278 -71 -262 -37
rect -328 -87 -262 -71
rect -210 -37 -144 -21
rect -210 -71 -194 -37
rect -160 -71 -144 -37
rect -210 -87 -144 -71
rect -92 -37 -26 -21
rect -92 -71 -76 -37
rect -42 -71 -26 -37
rect -92 -87 -26 -71
rect 26 -37 92 -21
rect 26 -71 42 -37
rect 76 -71 92 -37
rect 26 -87 92 -71
rect 144 -37 210 -21
rect 144 -71 160 -37
rect 194 -71 210 -37
rect 144 -87 210 -71
rect 262 -37 328 -21
rect 262 -71 278 -37
rect 312 -71 328 -37
rect 262 -87 328 -71
rect 380 -37 446 -21
rect 380 -71 396 -37
rect 430 -71 446 -37
rect 380 -87 446 -71
rect 498 -37 564 -21
rect 498 -71 514 -37
rect 548 -71 564 -37
rect 498 -87 564 -71
rect 616 -37 682 -21
rect 616 -71 632 -37
rect 666 -71 682 -37
rect 616 -87 682 -71
rect 734 -37 800 -21
rect 734 -71 750 -37
rect 784 -71 800 -37
rect 734 -87 800 -71
rect 852 -37 918 -21
rect 852 -71 868 -37
rect 902 -71 918 -37
rect 852 -87 918 -71
rect 970 -37 1036 -21
rect 970 -71 986 -37
rect 1020 -71 1036 -37
rect 970 -87 1036 -71
rect 1088 -37 1154 -21
rect 1088 -71 1104 -37
rect 1138 -71 1154 -37
rect 1088 -87 1154 -71
rect 1206 -37 1272 -21
rect 1206 -71 1222 -37
rect 1256 -71 1272 -37
rect 1206 -87 1272 -71
rect 1324 -37 1390 -21
rect 1324 -71 1340 -37
rect 1374 -71 1390 -37
rect 1324 -87 1390 -71
rect 1442 -37 1508 -21
rect 1442 -71 1458 -37
rect 1492 -71 1508 -37
rect 1442 -87 1508 -71
rect 1560 -37 1626 -21
rect 1560 -71 1576 -37
rect 1610 -71 1626 -37
rect 1560 -87 1626 -71
rect 1678 -37 1744 -21
rect 1678 -71 1694 -37
rect 1728 -71 1744 -37
rect 1678 -87 1744 -71
rect 1796 -37 1862 -21
rect 1796 -71 1812 -37
rect 1846 -71 1862 -37
rect 1796 -87 1862 -71
rect 1914 -37 1980 -21
rect 1914 -71 1930 -37
rect 1964 -71 1980 -37
rect 1914 -87 1980 -71
rect 2032 -37 2098 -21
rect 2032 -71 2048 -37
rect 2082 -71 2098 -37
rect 2032 -87 2098 -71
rect 2150 -37 2216 -21
rect 2150 -71 2166 -37
rect 2200 -71 2216 -37
rect 2150 -87 2216 -71
rect 2268 -37 2334 -21
rect 2268 -71 2284 -37
rect 2318 -71 2334 -37
rect 2268 -87 2334 -71
rect 2386 -37 2452 -21
rect 2386 -71 2402 -37
rect 2436 -71 2452 -37
rect 2386 -87 2452 -71
rect 2504 -37 2570 -21
rect 2504 -71 2520 -37
rect 2554 -71 2570 -37
rect 2504 -87 2570 -71
rect 2622 -37 2688 -21
rect 2622 -71 2638 -37
rect 2672 -71 2688 -37
rect 2622 -87 2688 -71
rect 2740 -37 2806 -21
rect 2740 -71 2756 -37
rect 2790 -71 2806 -37
rect 2740 -87 2806 -71
rect 2858 -37 2924 -21
rect 2858 -71 2874 -37
rect 2908 -71 2924 -37
rect 2858 -87 2924 -71
rect -2921 -118 -2861 -87
rect -2803 -118 -2743 -87
rect -2685 -118 -2625 -87
rect -2567 -118 -2507 -87
rect -2449 -118 -2389 -87
rect -2331 -118 -2271 -87
rect -2213 -118 -2153 -87
rect -2095 -118 -2035 -87
rect -1977 -118 -1917 -87
rect -1859 -118 -1799 -87
rect -1741 -118 -1681 -87
rect -1623 -118 -1563 -87
rect -1505 -118 -1445 -87
rect -1387 -118 -1327 -87
rect -1269 -118 -1209 -87
rect -1151 -118 -1091 -87
rect -1033 -118 -973 -87
rect -915 -118 -855 -87
rect -797 -118 -737 -87
rect -679 -118 -619 -87
rect -561 -118 -501 -87
rect -443 -118 -383 -87
rect -325 -118 -265 -87
rect -207 -118 -147 -87
rect -89 -118 -29 -87
rect 29 -118 89 -87
rect 147 -118 207 -87
rect 265 -118 325 -87
rect 383 -118 443 -87
rect 501 -118 561 -87
rect 619 -118 679 -87
rect 737 -118 797 -87
rect 855 -118 915 -87
rect 973 -118 1033 -87
rect 1091 -118 1151 -87
rect 1209 -118 1269 -87
rect 1327 -118 1387 -87
rect 1445 -118 1505 -87
rect 1563 -118 1623 -87
rect 1681 -118 1741 -87
rect 1799 -118 1859 -87
rect 1917 -118 1977 -87
rect 2035 -118 2095 -87
rect 2153 -118 2213 -87
rect 2271 -118 2331 -87
rect 2389 -118 2449 -87
rect 2507 -118 2567 -87
rect 2625 -118 2685 -87
rect 2743 -118 2803 -87
rect 2861 -118 2921 -87
rect -2921 -749 -2861 -718
rect -2803 -749 -2743 -718
rect -2685 -749 -2625 -718
rect -2567 -749 -2507 -718
rect -2449 -749 -2389 -718
rect -2331 -749 -2271 -718
rect -2213 -749 -2153 -718
rect -2095 -749 -2035 -718
rect -1977 -749 -1917 -718
rect -1859 -749 -1799 -718
rect -1741 -749 -1681 -718
rect -1623 -749 -1563 -718
rect -1505 -749 -1445 -718
rect -1387 -749 -1327 -718
rect -1269 -749 -1209 -718
rect -1151 -749 -1091 -718
rect -1033 -749 -973 -718
rect -915 -749 -855 -718
rect -797 -749 -737 -718
rect -679 -749 -619 -718
rect -561 -749 -501 -718
rect -443 -749 -383 -718
rect -325 -749 -265 -718
rect -207 -749 -147 -718
rect -89 -749 -29 -718
rect 29 -749 89 -718
rect 147 -749 207 -718
rect 265 -749 325 -718
rect 383 -749 443 -718
rect 501 -749 561 -718
rect 619 -749 679 -718
rect 737 -749 797 -718
rect 855 -749 915 -718
rect 973 -749 1033 -718
rect 1091 -749 1151 -718
rect 1209 -749 1269 -718
rect 1327 -749 1387 -718
rect 1445 -749 1505 -718
rect 1563 -749 1623 -718
rect 1681 -749 1741 -718
rect 1799 -749 1859 -718
rect 1917 -749 1977 -718
rect 2035 -749 2095 -718
rect 2153 -749 2213 -718
rect 2271 -749 2331 -718
rect 2389 -749 2449 -718
rect 2507 -749 2567 -718
rect 2625 -749 2685 -718
rect 2743 -749 2803 -718
rect 2861 -749 2921 -718
rect -2924 -765 -2858 -749
rect -2924 -799 -2908 -765
rect -2874 -799 -2858 -765
rect -2924 -815 -2858 -799
rect -2806 -765 -2740 -749
rect -2806 -799 -2790 -765
rect -2756 -799 -2740 -765
rect -2806 -815 -2740 -799
rect -2688 -765 -2622 -749
rect -2688 -799 -2672 -765
rect -2638 -799 -2622 -765
rect -2688 -815 -2622 -799
rect -2570 -765 -2504 -749
rect -2570 -799 -2554 -765
rect -2520 -799 -2504 -765
rect -2570 -815 -2504 -799
rect -2452 -765 -2386 -749
rect -2452 -799 -2436 -765
rect -2402 -799 -2386 -765
rect -2452 -815 -2386 -799
rect -2334 -765 -2268 -749
rect -2334 -799 -2318 -765
rect -2284 -799 -2268 -765
rect -2334 -815 -2268 -799
rect -2216 -765 -2150 -749
rect -2216 -799 -2200 -765
rect -2166 -799 -2150 -765
rect -2216 -815 -2150 -799
rect -2098 -765 -2032 -749
rect -2098 -799 -2082 -765
rect -2048 -799 -2032 -765
rect -2098 -815 -2032 -799
rect -1980 -765 -1914 -749
rect -1980 -799 -1964 -765
rect -1930 -799 -1914 -765
rect -1980 -815 -1914 -799
rect -1862 -765 -1796 -749
rect -1862 -799 -1846 -765
rect -1812 -799 -1796 -765
rect -1862 -815 -1796 -799
rect -1744 -765 -1678 -749
rect -1744 -799 -1728 -765
rect -1694 -799 -1678 -765
rect -1744 -815 -1678 -799
rect -1626 -765 -1560 -749
rect -1626 -799 -1610 -765
rect -1576 -799 -1560 -765
rect -1626 -815 -1560 -799
rect -1508 -765 -1442 -749
rect -1508 -799 -1492 -765
rect -1458 -799 -1442 -765
rect -1508 -815 -1442 -799
rect -1390 -765 -1324 -749
rect -1390 -799 -1374 -765
rect -1340 -799 -1324 -765
rect -1390 -815 -1324 -799
rect -1272 -765 -1206 -749
rect -1272 -799 -1256 -765
rect -1222 -799 -1206 -765
rect -1272 -815 -1206 -799
rect -1154 -765 -1088 -749
rect -1154 -799 -1138 -765
rect -1104 -799 -1088 -765
rect -1154 -815 -1088 -799
rect -1036 -765 -970 -749
rect -1036 -799 -1020 -765
rect -986 -799 -970 -765
rect -1036 -815 -970 -799
rect -918 -765 -852 -749
rect -918 -799 -902 -765
rect -868 -799 -852 -765
rect -918 -815 -852 -799
rect -800 -765 -734 -749
rect -800 -799 -784 -765
rect -750 -799 -734 -765
rect -800 -815 -734 -799
rect -682 -765 -616 -749
rect -682 -799 -666 -765
rect -632 -799 -616 -765
rect -682 -815 -616 -799
rect -564 -765 -498 -749
rect -564 -799 -548 -765
rect -514 -799 -498 -765
rect -564 -815 -498 -799
rect -446 -765 -380 -749
rect -446 -799 -430 -765
rect -396 -799 -380 -765
rect -446 -815 -380 -799
rect -328 -765 -262 -749
rect -328 -799 -312 -765
rect -278 -799 -262 -765
rect -328 -815 -262 -799
rect -210 -765 -144 -749
rect -210 -799 -194 -765
rect -160 -799 -144 -765
rect -210 -815 -144 -799
rect -92 -765 -26 -749
rect -92 -799 -76 -765
rect -42 -799 -26 -765
rect -92 -815 -26 -799
rect 26 -765 92 -749
rect 26 -799 42 -765
rect 76 -799 92 -765
rect 26 -815 92 -799
rect 144 -765 210 -749
rect 144 -799 160 -765
rect 194 -799 210 -765
rect 144 -815 210 -799
rect 262 -765 328 -749
rect 262 -799 278 -765
rect 312 -799 328 -765
rect 262 -815 328 -799
rect 380 -765 446 -749
rect 380 -799 396 -765
rect 430 -799 446 -765
rect 380 -815 446 -799
rect 498 -765 564 -749
rect 498 -799 514 -765
rect 548 -799 564 -765
rect 498 -815 564 -799
rect 616 -765 682 -749
rect 616 -799 632 -765
rect 666 -799 682 -765
rect 616 -815 682 -799
rect 734 -765 800 -749
rect 734 -799 750 -765
rect 784 -799 800 -765
rect 734 -815 800 -799
rect 852 -765 918 -749
rect 852 -799 868 -765
rect 902 -799 918 -765
rect 852 -815 918 -799
rect 970 -765 1036 -749
rect 970 -799 986 -765
rect 1020 -799 1036 -765
rect 970 -815 1036 -799
rect 1088 -765 1154 -749
rect 1088 -799 1104 -765
rect 1138 -799 1154 -765
rect 1088 -815 1154 -799
rect 1206 -765 1272 -749
rect 1206 -799 1222 -765
rect 1256 -799 1272 -765
rect 1206 -815 1272 -799
rect 1324 -765 1390 -749
rect 1324 -799 1340 -765
rect 1374 -799 1390 -765
rect 1324 -815 1390 -799
rect 1442 -765 1508 -749
rect 1442 -799 1458 -765
rect 1492 -799 1508 -765
rect 1442 -815 1508 -799
rect 1560 -765 1626 -749
rect 1560 -799 1576 -765
rect 1610 -799 1626 -765
rect 1560 -815 1626 -799
rect 1678 -765 1744 -749
rect 1678 -799 1694 -765
rect 1728 -799 1744 -765
rect 1678 -815 1744 -799
rect 1796 -765 1862 -749
rect 1796 -799 1812 -765
rect 1846 -799 1862 -765
rect 1796 -815 1862 -799
rect 1914 -765 1980 -749
rect 1914 -799 1930 -765
rect 1964 -799 1980 -765
rect 1914 -815 1980 -799
rect 2032 -765 2098 -749
rect 2032 -799 2048 -765
rect 2082 -799 2098 -765
rect 2032 -815 2098 -799
rect 2150 -765 2216 -749
rect 2150 -799 2166 -765
rect 2200 -799 2216 -765
rect 2150 -815 2216 -799
rect 2268 -765 2334 -749
rect 2268 -799 2284 -765
rect 2318 -799 2334 -765
rect 2268 -815 2334 -799
rect 2386 -765 2452 -749
rect 2386 -799 2402 -765
rect 2436 -799 2452 -765
rect 2386 -815 2452 -799
rect 2504 -765 2570 -749
rect 2504 -799 2520 -765
rect 2554 -799 2570 -765
rect 2504 -815 2570 -799
rect 2622 -765 2688 -749
rect 2622 -799 2638 -765
rect 2672 -799 2688 -765
rect 2622 -815 2688 -799
rect 2740 -765 2806 -749
rect 2740 -799 2756 -765
rect 2790 -799 2806 -765
rect 2740 -815 2806 -799
rect 2858 -765 2924 -749
rect 2858 -799 2874 -765
rect 2908 -799 2924 -765
rect 2858 -815 2924 -799
rect -2924 -873 -2858 -857
rect -2924 -907 -2908 -873
rect -2874 -907 -2858 -873
rect -2924 -923 -2858 -907
rect -2806 -873 -2740 -857
rect -2806 -907 -2790 -873
rect -2756 -907 -2740 -873
rect -2806 -923 -2740 -907
rect -2688 -873 -2622 -857
rect -2688 -907 -2672 -873
rect -2638 -907 -2622 -873
rect -2688 -923 -2622 -907
rect -2570 -873 -2504 -857
rect -2570 -907 -2554 -873
rect -2520 -907 -2504 -873
rect -2570 -923 -2504 -907
rect -2452 -873 -2386 -857
rect -2452 -907 -2436 -873
rect -2402 -907 -2386 -873
rect -2452 -923 -2386 -907
rect -2334 -873 -2268 -857
rect -2334 -907 -2318 -873
rect -2284 -907 -2268 -873
rect -2334 -923 -2268 -907
rect -2216 -873 -2150 -857
rect -2216 -907 -2200 -873
rect -2166 -907 -2150 -873
rect -2216 -923 -2150 -907
rect -2098 -873 -2032 -857
rect -2098 -907 -2082 -873
rect -2048 -907 -2032 -873
rect -2098 -923 -2032 -907
rect -1980 -873 -1914 -857
rect -1980 -907 -1964 -873
rect -1930 -907 -1914 -873
rect -1980 -923 -1914 -907
rect -1862 -873 -1796 -857
rect -1862 -907 -1846 -873
rect -1812 -907 -1796 -873
rect -1862 -923 -1796 -907
rect -1744 -873 -1678 -857
rect -1744 -907 -1728 -873
rect -1694 -907 -1678 -873
rect -1744 -923 -1678 -907
rect -1626 -873 -1560 -857
rect -1626 -907 -1610 -873
rect -1576 -907 -1560 -873
rect -1626 -923 -1560 -907
rect -1508 -873 -1442 -857
rect -1508 -907 -1492 -873
rect -1458 -907 -1442 -873
rect -1508 -923 -1442 -907
rect -1390 -873 -1324 -857
rect -1390 -907 -1374 -873
rect -1340 -907 -1324 -873
rect -1390 -923 -1324 -907
rect -1272 -873 -1206 -857
rect -1272 -907 -1256 -873
rect -1222 -907 -1206 -873
rect -1272 -923 -1206 -907
rect -1154 -873 -1088 -857
rect -1154 -907 -1138 -873
rect -1104 -907 -1088 -873
rect -1154 -923 -1088 -907
rect -1036 -873 -970 -857
rect -1036 -907 -1020 -873
rect -986 -907 -970 -873
rect -1036 -923 -970 -907
rect -918 -873 -852 -857
rect -918 -907 -902 -873
rect -868 -907 -852 -873
rect -918 -923 -852 -907
rect -800 -873 -734 -857
rect -800 -907 -784 -873
rect -750 -907 -734 -873
rect -800 -923 -734 -907
rect -682 -873 -616 -857
rect -682 -907 -666 -873
rect -632 -907 -616 -873
rect -682 -923 -616 -907
rect -564 -873 -498 -857
rect -564 -907 -548 -873
rect -514 -907 -498 -873
rect -564 -923 -498 -907
rect -446 -873 -380 -857
rect -446 -907 -430 -873
rect -396 -907 -380 -873
rect -446 -923 -380 -907
rect -328 -873 -262 -857
rect -328 -907 -312 -873
rect -278 -907 -262 -873
rect -328 -923 -262 -907
rect -210 -873 -144 -857
rect -210 -907 -194 -873
rect -160 -907 -144 -873
rect -210 -923 -144 -907
rect -92 -873 -26 -857
rect -92 -907 -76 -873
rect -42 -907 -26 -873
rect -92 -923 -26 -907
rect 26 -873 92 -857
rect 26 -907 42 -873
rect 76 -907 92 -873
rect 26 -923 92 -907
rect 144 -873 210 -857
rect 144 -907 160 -873
rect 194 -907 210 -873
rect 144 -923 210 -907
rect 262 -873 328 -857
rect 262 -907 278 -873
rect 312 -907 328 -873
rect 262 -923 328 -907
rect 380 -873 446 -857
rect 380 -907 396 -873
rect 430 -907 446 -873
rect 380 -923 446 -907
rect 498 -873 564 -857
rect 498 -907 514 -873
rect 548 -907 564 -873
rect 498 -923 564 -907
rect 616 -873 682 -857
rect 616 -907 632 -873
rect 666 -907 682 -873
rect 616 -923 682 -907
rect 734 -873 800 -857
rect 734 -907 750 -873
rect 784 -907 800 -873
rect 734 -923 800 -907
rect 852 -873 918 -857
rect 852 -907 868 -873
rect 902 -907 918 -873
rect 852 -923 918 -907
rect 970 -873 1036 -857
rect 970 -907 986 -873
rect 1020 -907 1036 -873
rect 970 -923 1036 -907
rect 1088 -873 1154 -857
rect 1088 -907 1104 -873
rect 1138 -907 1154 -873
rect 1088 -923 1154 -907
rect 1206 -873 1272 -857
rect 1206 -907 1222 -873
rect 1256 -907 1272 -873
rect 1206 -923 1272 -907
rect 1324 -873 1390 -857
rect 1324 -907 1340 -873
rect 1374 -907 1390 -873
rect 1324 -923 1390 -907
rect 1442 -873 1508 -857
rect 1442 -907 1458 -873
rect 1492 -907 1508 -873
rect 1442 -923 1508 -907
rect 1560 -873 1626 -857
rect 1560 -907 1576 -873
rect 1610 -907 1626 -873
rect 1560 -923 1626 -907
rect 1678 -873 1744 -857
rect 1678 -907 1694 -873
rect 1728 -907 1744 -873
rect 1678 -923 1744 -907
rect 1796 -873 1862 -857
rect 1796 -907 1812 -873
rect 1846 -907 1862 -873
rect 1796 -923 1862 -907
rect 1914 -873 1980 -857
rect 1914 -907 1930 -873
rect 1964 -907 1980 -873
rect 1914 -923 1980 -907
rect 2032 -873 2098 -857
rect 2032 -907 2048 -873
rect 2082 -907 2098 -873
rect 2032 -923 2098 -907
rect 2150 -873 2216 -857
rect 2150 -907 2166 -873
rect 2200 -907 2216 -873
rect 2150 -923 2216 -907
rect 2268 -873 2334 -857
rect 2268 -907 2284 -873
rect 2318 -907 2334 -873
rect 2268 -923 2334 -907
rect 2386 -873 2452 -857
rect 2386 -907 2402 -873
rect 2436 -907 2452 -873
rect 2386 -923 2452 -907
rect 2504 -873 2570 -857
rect 2504 -907 2520 -873
rect 2554 -907 2570 -873
rect 2504 -923 2570 -907
rect 2622 -873 2688 -857
rect 2622 -907 2638 -873
rect 2672 -907 2688 -873
rect 2622 -923 2688 -907
rect 2740 -873 2806 -857
rect 2740 -907 2756 -873
rect 2790 -907 2806 -873
rect 2740 -923 2806 -907
rect 2858 -873 2924 -857
rect 2858 -907 2874 -873
rect 2908 -907 2924 -873
rect 2858 -923 2924 -907
rect -2921 -954 -2861 -923
rect -2803 -954 -2743 -923
rect -2685 -954 -2625 -923
rect -2567 -954 -2507 -923
rect -2449 -954 -2389 -923
rect -2331 -954 -2271 -923
rect -2213 -954 -2153 -923
rect -2095 -954 -2035 -923
rect -1977 -954 -1917 -923
rect -1859 -954 -1799 -923
rect -1741 -954 -1681 -923
rect -1623 -954 -1563 -923
rect -1505 -954 -1445 -923
rect -1387 -954 -1327 -923
rect -1269 -954 -1209 -923
rect -1151 -954 -1091 -923
rect -1033 -954 -973 -923
rect -915 -954 -855 -923
rect -797 -954 -737 -923
rect -679 -954 -619 -923
rect -561 -954 -501 -923
rect -443 -954 -383 -923
rect -325 -954 -265 -923
rect -207 -954 -147 -923
rect -89 -954 -29 -923
rect 29 -954 89 -923
rect 147 -954 207 -923
rect 265 -954 325 -923
rect 383 -954 443 -923
rect 501 -954 561 -923
rect 619 -954 679 -923
rect 737 -954 797 -923
rect 855 -954 915 -923
rect 973 -954 1033 -923
rect 1091 -954 1151 -923
rect 1209 -954 1269 -923
rect 1327 -954 1387 -923
rect 1445 -954 1505 -923
rect 1563 -954 1623 -923
rect 1681 -954 1741 -923
rect 1799 -954 1859 -923
rect 1917 -954 1977 -923
rect 2035 -954 2095 -923
rect 2153 -954 2213 -923
rect 2271 -954 2331 -923
rect 2389 -954 2449 -923
rect 2507 -954 2567 -923
rect 2625 -954 2685 -923
rect 2743 -954 2803 -923
rect 2861 -954 2921 -923
rect -2921 -1585 -2861 -1554
rect -2803 -1585 -2743 -1554
rect -2685 -1585 -2625 -1554
rect -2567 -1585 -2507 -1554
rect -2449 -1585 -2389 -1554
rect -2331 -1585 -2271 -1554
rect -2213 -1585 -2153 -1554
rect -2095 -1585 -2035 -1554
rect -1977 -1585 -1917 -1554
rect -1859 -1585 -1799 -1554
rect -1741 -1585 -1681 -1554
rect -1623 -1585 -1563 -1554
rect -1505 -1585 -1445 -1554
rect -1387 -1585 -1327 -1554
rect -1269 -1585 -1209 -1554
rect -1151 -1585 -1091 -1554
rect -1033 -1585 -973 -1554
rect -915 -1585 -855 -1554
rect -797 -1585 -737 -1554
rect -679 -1585 -619 -1554
rect -561 -1585 -501 -1554
rect -443 -1585 -383 -1554
rect -325 -1585 -265 -1554
rect -207 -1585 -147 -1554
rect -89 -1585 -29 -1554
rect 29 -1585 89 -1554
rect 147 -1585 207 -1554
rect 265 -1585 325 -1554
rect 383 -1585 443 -1554
rect 501 -1585 561 -1554
rect 619 -1585 679 -1554
rect 737 -1585 797 -1554
rect 855 -1585 915 -1554
rect 973 -1585 1033 -1554
rect 1091 -1585 1151 -1554
rect 1209 -1585 1269 -1554
rect 1327 -1585 1387 -1554
rect 1445 -1585 1505 -1554
rect 1563 -1585 1623 -1554
rect 1681 -1585 1741 -1554
rect 1799 -1585 1859 -1554
rect 1917 -1585 1977 -1554
rect 2035 -1585 2095 -1554
rect 2153 -1585 2213 -1554
rect 2271 -1585 2331 -1554
rect 2389 -1585 2449 -1554
rect 2507 -1585 2567 -1554
rect 2625 -1585 2685 -1554
rect 2743 -1585 2803 -1554
rect 2861 -1585 2921 -1554
rect -2924 -1601 -2858 -1585
rect -2924 -1635 -2908 -1601
rect -2874 -1635 -2858 -1601
rect -2924 -1651 -2858 -1635
rect -2806 -1601 -2740 -1585
rect -2806 -1635 -2790 -1601
rect -2756 -1635 -2740 -1601
rect -2806 -1651 -2740 -1635
rect -2688 -1601 -2622 -1585
rect -2688 -1635 -2672 -1601
rect -2638 -1635 -2622 -1601
rect -2688 -1651 -2622 -1635
rect -2570 -1601 -2504 -1585
rect -2570 -1635 -2554 -1601
rect -2520 -1635 -2504 -1601
rect -2570 -1651 -2504 -1635
rect -2452 -1601 -2386 -1585
rect -2452 -1635 -2436 -1601
rect -2402 -1635 -2386 -1601
rect -2452 -1651 -2386 -1635
rect -2334 -1601 -2268 -1585
rect -2334 -1635 -2318 -1601
rect -2284 -1635 -2268 -1601
rect -2334 -1651 -2268 -1635
rect -2216 -1601 -2150 -1585
rect -2216 -1635 -2200 -1601
rect -2166 -1635 -2150 -1601
rect -2216 -1651 -2150 -1635
rect -2098 -1601 -2032 -1585
rect -2098 -1635 -2082 -1601
rect -2048 -1635 -2032 -1601
rect -2098 -1651 -2032 -1635
rect -1980 -1601 -1914 -1585
rect -1980 -1635 -1964 -1601
rect -1930 -1635 -1914 -1601
rect -1980 -1651 -1914 -1635
rect -1862 -1601 -1796 -1585
rect -1862 -1635 -1846 -1601
rect -1812 -1635 -1796 -1601
rect -1862 -1651 -1796 -1635
rect -1744 -1601 -1678 -1585
rect -1744 -1635 -1728 -1601
rect -1694 -1635 -1678 -1601
rect -1744 -1651 -1678 -1635
rect -1626 -1601 -1560 -1585
rect -1626 -1635 -1610 -1601
rect -1576 -1635 -1560 -1601
rect -1626 -1651 -1560 -1635
rect -1508 -1601 -1442 -1585
rect -1508 -1635 -1492 -1601
rect -1458 -1635 -1442 -1601
rect -1508 -1651 -1442 -1635
rect -1390 -1601 -1324 -1585
rect -1390 -1635 -1374 -1601
rect -1340 -1635 -1324 -1601
rect -1390 -1651 -1324 -1635
rect -1272 -1601 -1206 -1585
rect -1272 -1635 -1256 -1601
rect -1222 -1635 -1206 -1601
rect -1272 -1651 -1206 -1635
rect -1154 -1601 -1088 -1585
rect -1154 -1635 -1138 -1601
rect -1104 -1635 -1088 -1601
rect -1154 -1651 -1088 -1635
rect -1036 -1601 -970 -1585
rect -1036 -1635 -1020 -1601
rect -986 -1635 -970 -1601
rect -1036 -1651 -970 -1635
rect -918 -1601 -852 -1585
rect -918 -1635 -902 -1601
rect -868 -1635 -852 -1601
rect -918 -1651 -852 -1635
rect -800 -1601 -734 -1585
rect -800 -1635 -784 -1601
rect -750 -1635 -734 -1601
rect -800 -1651 -734 -1635
rect -682 -1601 -616 -1585
rect -682 -1635 -666 -1601
rect -632 -1635 -616 -1601
rect -682 -1651 -616 -1635
rect -564 -1601 -498 -1585
rect -564 -1635 -548 -1601
rect -514 -1635 -498 -1601
rect -564 -1651 -498 -1635
rect -446 -1601 -380 -1585
rect -446 -1635 -430 -1601
rect -396 -1635 -380 -1601
rect -446 -1651 -380 -1635
rect -328 -1601 -262 -1585
rect -328 -1635 -312 -1601
rect -278 -1635 -262 -1601
rect -328 -1651 -262 -1635
rect -210 -1601 -144 -1585
rect -210 -1635 -194 -1601
rect -160 -1635 -144 -1601
rect -210 -1651 -144 -1635
rect -92 -1601 -26 -1585
rect -92 -1635 -76 -1601
rect -42 -1635 -26 -1601
rect -92 -1651 -26 -1635
rect 26 -1601 92 -1585
rect 26 -1635 42 -1601
rect 76 -1635 92 -1601
rect 26 -1651 92 -1635
rect 144 -1601 210 -1585
rect 144 -1635 160 -1601
rect 194 -1635 210 -1601
rect 144 -1651 210 -1635
rect 262 -1601 328 -1585
rect 262 -1635 278 -1601
rect 312 -1635 328 -1601
rect 262 -1651 328 -1635
rect 380 -1601 446 -1585
rect 380 -1635 396 -1601
rect 430 -1635 446 -1601
rect 380 -1651 446 -1635
rect 498 -1601 564 -1585
rect 498 -1635 514 -1601
rect 548 -1635 564 -1601
rect 498 -1651 564 -1635
rect 616 -1601 682 -1585
rect 616 -1635 632 -1601
rect 666 -1635 682 -1601
rect 616 -1651 682 -1635
rect 734 -1601 800 -1585
rect 734 -1635 750 -1601
rect 784 -1635 800 -1601
rect 734 -1651 800 -1635
rect 852 -1601 918 -1585
rect 852 -1635 868 -1601
rect 902 -1635 918 -1601
rect 852 -1651 918 -1635
rect 970 -1601 1036 -1585
rect 970 -1635 986 -1601
rect 1020 -1635 1036 -1601
rect 970 -1651 1036 -1635
rect 1088 -1601 1154 -1585
rect 1088 -1635 1104 -1601
rect 1138 -1635 1154 -1601
rect 1088 -1651 1154 -1635
rect 1206 -1601 1272 -1585
rect 1206 -1635 1222 -1601
rect 1256 -1635 1272 -1601
rect 1206 -1651 1272 -1635
rect 1324 -1601 1390 -1585
rect 1324 -1635 1340 -1601
rect 1374 -1635 1390 -1601
rect 1324 -1651 1390 -1635
rect 1442 -1601 1508 -1585
rect 1442 -1635 1458 -1601
rect 1492 -1635 1508 -1601
rect 1442 -1651 1508 -1635
rect 1560 -1601 1626 -1585
rect 1560 -1635 1576 -1601
rect 1610 -1635 1626 -1601
rect 1560 -1651 1626 -1635
rect 1678 -1601 1744 -1585
rect 1678 -1635 1694 -1601
rect 1728 -1635 1744 -1601
rect 1678 -1651 1744 -1635
rect 1796 -1601 1862 -1585
rect 1796 -1635 1812 -1601
rect 1846 -1635 1862 -1601
rect 1796 -1651 1862 -1635
rect 1914 -1601 1980 -1585
rect 1914 -1635 1930 -1601
rect 1964 -1635 1980 -1601
rect 1914 -1651 1980 -1635
rect 2032 -1601 2098 -1585
rect 2032 -1635 2048 -1601
rect 2082 -1635 2098 -1601
rect 2032 -1651 2098 -1635
rect 2150 -1601 2216 -1585
rect 2150 -1635 2166 -1601
rect 2200 -1635 2216 -1601
rect 2150 -1651 2216 -1635
rect 2268 -1601 2334 -1585
rect 2268 -1635 2284 -1601
rect 2318 -1635 2334 -1601
rect 2268 -1651 2334 -1635
rect 2386 -1601 2452 -1585
rect 2386 -1635 2402 -1601
rect 2436 -1635 2452 -1601
rect 2386 -1651 2452 -1635
rect 2504 -1601 2570 -1585
rect 2504 -1635 2520 -1601
rect 2554 -1635 2570 -1601
rect 2504 -1651 2570 -1635
rect 2622 -1601 2688 -1585
rect 2622 -1635 2638 -1601
rect 2672 -1635 2688 -1601
rect 2622 -1651 2688 -1635
rect 2740 -1601 2806 -1585
rect 2740 -1635 2756 -1601
rect 2790 -1635 2806 -1601
rect 2740 -1651 2806 -1635
rect 2858 -1601 2924 -1585
rect 2858 -1635 2874 -1601
rect 2908 -1635 2924 -1601
rect 2858 -1651 2924 -1635
<< polycont >>
rect -2908 1601 -2874 1635
rect -2790 1601 -2756 1635
rect -2672 1601 -2638 1635
rect -2554 1601 -2520 1635
rect -2436 1601 -2402 1635
rect -2318 1601 -2284 1635
rect -2200 1601 -2166 1635
rect -2082 1601 -2048 1635
rect -1964 1601 -1930 1635
rect -1846 1601 -1812 1635
rect -1728 1601 -1694 1635
rect -1610 1601 -1576 1635
rect -1492 1601 -1458 1635
rect -1374 1601 -1340 1635
rect -1256 1601 -1222 1635
rect -1138 1601 -1104 1635
rect -1020 1601 -986 1635
rect -902 1601 -868 1635
rect -784 1601 -750 1635
rect -666 1601 -632 1635
rect -548 1601 -514 1635
rect -430 1601 -396 1635
rect -312 1601 -278 1635
rect -194 1601 -160 1635
rect -76 1601 -42 1635
rect 42 1601 76 1635
rect 160 1601 194 1635
rect 278 1601 312 1635
rect 396 1601 430 1635
rect 514 1601 548 1635
rect 632 1601 666 1635
rect 750 1601 784 1635
rect 868 1601 902 1635
rect 986 1601 1020 1635
rect 1104 1601 1138 1635
rect 1222 1601 1256 1635
rect 1340 1601 1374 1635
rect 1458 1601 1492 1635
rect 1576 1601 1610 1635
rect 1694 1601 1728 1635
rect 1812 1601 1846 1635
rect 1930 1601 1964 1635
rect 2048 1601 2082 1635
rect 2166 1601 2200 1635
rect 2284 1601 2318 1635
rect 2402 1601 2436 1635
rect 2520 1601 2554 1635
rect 2638 1601 2672 1635
rect 2756 1601 2790 1635
rect 2874 1601 2908 1635
rect -2908 873 -2874 907
rect -2790 873 -2756 907
rect -2672 873 -2638 907
rect -2554 873 -2520 907
rect -2436 873 -2402 907
rect -2318 873 -2284 907
rect -2200 873 -2166 907
rect -2082 873 -2048 907
rect -1964 873 -1930 907
rect -1846 873 -1812 907
rect -1728 873 -1694 907
rect -1610 873 -1576 907
rect -1492 873 -1458 907
rect -1374 873 -1340 907
rect -1256 873 -1222 907
rect -1138 873 -1104 907
rect -1020 873 -986 907
rect -902 873 -868 907
rect -784 873 -750 907
rect -666 873 -632 907
rect -548 873 -514 907
rect -430 873 -396 907
rect -312 873 -278 907
rect -194 873 -160 907
rect -76 873 -42 907
rect 42 873 76 907
rect 160 873 194 907
rect 278 873 312 907
rect 396 873 430 907
rect 514 873 548 907
rect 632 873 666 907
rect 750 873 784 907
rect 868 873 902 907
rect 986 873 1020 907
rect 1104 873 1138 907
rect 1222 873 1256 907
rect 1340 873 1374 907
rect 1458 873 1492 907
rect 1576 873 1610 907
rect 1694 873 1728 907
rect 1812 873 1846 907
rect 1930 873 1964 907
rect 2048 873 2082 907
rect 2166 873 2200 907
rect 2284 873 2318 907
rect 2402 873 2436 907
rect 2520 873 2554 907
rect 2638 873 2672 907
rect 2756 873 2790 907
rect 2874 873 2908 907
rect -2908 765 -2874 799
rect -2790 765 -2756 799
rect -2672 765 -2638 799
rect -2554 765 -2520 799
rect -2436 765 -2402 799
rect -2318 765 -2284 799
rect -2200 765 -2166 799
rect -2082 765 -2048 799
rect -1964 765 -1930 799
rect -1846 765 -1812 799
rect -1728 765 -1694 799
rect -1610 765 -1576 799
rect -1492 765 -1458 799
rect -1374 765 -1340 799
rect -1256 765 -1222 799
rect -1138 765 -1104 799
rect -1020 765 -986 799
rect -902 765 -868 799
rect -784 765 -750 799
rect -666 765 -632 799
rect -548 765 -514 799
rect -430 765 -396 799
rect -312 765 -278 799
rect -194 765 -160 799
rect -76 765 -42 799
rect 42 765 76 799
rect 160 765 194 799
rect 278 765 312 799
rect 396 765 430 799
rect 514 765 548 799
rect 632 765 666 799
rect 750 765 784 799
rect 868 765 902 799
rect 986 765 1020 799
rect 1104 765 1138 799
rect 1222 765 1256 799
rect 1340 765 1374 799
rect 1458 765 1492 799
rect 1576 765 1610 799
rect 1694 765 1728 799
rect 1812 765 1846 799
rect 1930 765 1964 799
rect 2048 765 2082 799
rect 2166 765 2200 799
rect 2284 765 2318 799
rect 2402 765 2436 799
rect 2520 765 2554 799
rect 2638 765 2672 799
rect 2756 765 2790 799
rect 2874 765 2908 799
rect -2908 37 -2874 71
rect -2790 37 -2756 71
rect -2672 37 -2638 71
rect -2554 37 -2520 71
rect -2436 37 -2402 71
rect -2318 37 -2284 71
rect -2200 37 -2166 71
rect -2082 37 -2048 71
rect -1964 37 -1930 71
rect -1846 37 -1812 71
rect -1728 37 -1694 71
rect -1610 37 -1576 71
rect -1492 37 -1458 71
rect -1374 37 -1340 71
rect -1256 37 -1222 71
rect -1138 37 -1104 71
rect -1020 37 -986 71
rect -902 37 -868 71
rect -784 37 -750 71
rect -666 37 -632 71
rect -548 37 -514 71
rect -430 37 -396 71
rect -312 37 -278 71
rect -194 37 -160 71
rect -76 37 -42 71
rect 42 37 76 71
rect 160 37 194 71
rect 278 37 312 71
rect 396 37 430 71
rect 514 37 548 71
rect 632 37 666 71
rect 750 37 784 71
rect 868 37 902 71
rect 986 37 1020 71
rect 1104 37 1138 71
rect 1222 37 1256 71
rect 1340 37 1374 71
rect 1458 37 1492 71
rect 1576 37 1610 71
rect 1694 37 1728 71
rect 1812 37 1846 71
rect 1930 37 1964 71
rect 2048 37 2082 71
rect 2166 37 2200 71
rect 2284 37 2318 71
rect 2402 37 2436 71
rect 2520 37 2554 71
rect 2638 37 2672 71
rect 2756 37 2790 71
rect 2874 37 2908 71
rect -2908 -71 -2874 -37
rect -2790 -71 -2756 -37
rect -2672 -71 -2638 -37
rect -2554 -71 -2520 -37
rect -2436 -71 -2402 -37
rect -2318 -71 -2284 -37
rect -2200 -71 -2166 -37
rect -2082 -71 -2048 -37
rect -1964 -71 -1930 -37
rect -1846 -71 -1812 -37
rect -1728 -71 -1694 -37
rect -1610 -71 -1576 -37
rect -1492 -71 -1458 -37
rect -1374 -71 -1340 -37
rect -1256 -71 -1222 -37
rect -1138 -71 -1104 -37
rect -1020 -71 -986 -37
rect -902 -71 -868 -37
rect -784 -71 -750 -37
rect -666 -71 -632 -37
rect -548 -71 -514 -37
rect -430 -71 -396 -37
rect -312 -71 -278 -37
rect -194 -71 -160 -37
rect -76 -71 -42 -37
rect 42 -71 76 -37
rect 160 -71 194 -37
rect 278 -71 312 -37
rect 396 -71 430 -37
rect 514 -71 548 -37
rect 632 -71 666 -37
rect 750 -71 784 -37
rect 868 -71 902 -37
rect 986 -71 1020 -37
rect 1104 -71 1138 -37
rect 1222 -71 1256 -37
rect 1340 -71 1374 -37
rect 1458 -71 1492 -37
rect 1576 -71 1610 -37
rect 1694 -71 1728 -37
rect 1812 -71 1846 -37
rect 1930 -71 1964 -37
rect 2048 -71 2082 -37
rect 2166 -71 2200 -37
rect 2284 -71 2318 -37
rect 2402 -71 2436 -37
rect 2520 -71 2554 -37
rect 2638 -71 2672 -37
rect 2756 -71 2790 -37
rect 2874 -71 2908 -37
rect -2908 -799 -2874 -765
rect -2790 -799 -2756 -765
rect -2672 -799 -2638 -765
rect -2554 -799 -2520 -765
rect -2436 -799 -2402 -765
rect -2318 -799 -2284 -765
rect -2200 -799 -2166 -765
rect -2082 -799 -2048 -765
rect -1964 -799 -1930 -765
rect -1846 -799 -1812 -765
rect -1728 -799 -1694 -765
rect -1610 -799 -1576 -765
rect -1492 -799 -1458 -765
rect -1374 -799 -1340 -765
rect -1256 -799 -1222 -765
rect -1138 -799 -1104 -765
rect -1020 -799 -986 -765
rect -902 -799 -868 -765
rect -784 -799 -750 -765
rect -666 -799 -632 -765
rect -548 -799 -514 -765
rect -430 -799 -396 -765
rect -312 -799 -278 -765
rect -194 -799 -160 -765
rect -76 -799 -42 -765
rect 42 -799 76 -765
rect 160 -799 194 -765
rect 278 -799 312 -765
rect 396 -799 430 -765
rect 514 -799 548 -765
rect 632 -799 666 -765
rect 750 -799 784 -765
rect 868 -799 902 -765
rect 986 -799 1020 -765
rect 1104 -799 1138 -765
rect 1222 -799 1256 -765
rect 1340 -799 1374 -765
rect 1458 -799 1492 -765
rect 1576 -799 1610 -765
rect 1694 -799 1728 -765
rect 1812 -799 1846 -765
rect 1930 -799 1964 -765
rect 2048 -799 2082 -765
rect 2166 -799 2200 -765
rect 2284 -799 2318 -765
rect 2402 -799 2436 -765
rect 2520 -799 2554 -765
rect 2638 -799 2672 -765
rect 2756 -799 2790 -765
rect 2874 -799 2908 -765
rect -2908 -907 -2874 -873
rect -2790 -907 -2756 -873
rect -2672 -907 -2638 -873
rect -2554 -907 -2520 -873
rect -2436 -907 -2402 -873
rect -2318 -907 -2284 -873
rect -2200 -907 -2166 -873
rect -2082 -907 -2048 -873
rect -1964 -907 -1930 -873
rect -1846 -907 -1812 -873
rect -1728 -907 -1694 -873
rect -1610 -907 -1576 -873
rect -1492 -907 -1458 -873
rect -1374 -907 -1340 -873
rect -1256 -907 -1222 -873
rect -1138 -907 -1104 -873
rect -1020 -907 -986 -873
rect -902 -907 -868 -873
rect -784 -907 -750 -873
rect -666 -907 -632 -873
rect -548 -907 -514 -873
rect -430 -907 -396 -873
rect -312 -907 -278 -873
rect -194 -907 -160 -873
rect -76 -907 -42 -873
rect 42 -907 76 -873
rect 160 -907 194 -873
rect 278 -907 312 -873
rect 396 -907 430 -873
rect 514 -907 548 -873
rect 632 -907 666 -873
rect 750 -907 784 -873
rect 868 -907 902 -873
rect 986 -907 1020 -873
rect 1104 -907 1138 -873
rect 1222 -907 1256 -873
rect 1340 -907 1374 -873
rect 1458 -907 1492 -873
rect 1576 -907 1610 -873
rect 1694 -907 1728 -873
rect 1812 -907 1846 -873
rect 1930 -907 1964 -873
rect 2048 -907 2082 -873
rect 2166 -907 2200 -873
rect 2284 -907 2318 -873
rect 2402 -907 2436 -873
rect 2520 -907 2554 -873
rect 2638 -907 2672 -873
rect 2756 -907 2790 -873
rect 2874 -907 2908 -873
rect -2908 -1635 -2874 -1601
rect -2790 -1635 -2756 -1601
rect -2672 -1635 -2638 -1601
rect -2554 -1635 -2520 -1601
rect -2436 -1635 -2402 -1601
rect -2318 -1635 -2284 -1601
rect -2200 -1635 -2166 -1601
rect -2082 -1635 -2048 -1601
rect -1964 -1635 -1930 -1601
rect -1846 -1635 -1812 -1601
rect -1728 -1635 -1694 -1601
rect -1610 -1635 -1576 -1601
rect -1492 -1635 -1458 -1601
rect -1374 -1635 -1340 -1601
rect -1256 -1635 -1222 -1601
rect -1138 -1635 -1104 -1601
rect -1020 -1635 -986 -1601
rect -902 -1635 -868 -1601
rect -784 -1635 -750 -1601
rect -666 -1635 -632 -1601
rect -548 -1635 -514 -1601
rect -430 -1635 -396 -1601
rect -312 -1635 -278 -1601
rect -194 -1635 -160 -1601
rect -76 -1635 -42 -1601
rect 42 -1635 76 -1601
rect 160 -1635 194 -1601
rect 278 -1635 312 -1601
rect 396 -1635 430 -1601
rect 514 -1635 548 -1601
rect 632 -1635 666 -1601
rect 750 -1635 784 -1601
rect 868 -1635 902 -1601
rect 986 -1635 1020 -1601
rect 1104 -1635 1138 -1601
rect 1222 -1635 1256 -1601
rect 1340 -1635 1374 -1601
rect 1458 -1635 1492 -1601
rect 1576 -1635 1610 -1601
rect 1694 -1635 1728 -1601
rect 1812 -1635 1846 -1601
rect 1930 -1635 1964 -1601
rect 2048 -1635 2082 -1601
rect 2166 -1635 2200 -1601
rect 2284 -1635 2318 -1601
rect 2402 -1635 2436 -1601
rect 2520 -1635 2554 -1601
rect 2638 -1635 2672 -1601
rect 2756 -1635 2790 -1601
rect 2874 -1635 2908 -1601
<< locali >>
rect -3081 1703 -2985 1737
rect 2985 1703 3081 1737
rect -3081 1641 -3047 1703
rect 3047 1641 3081 1703
rect -2924 1601 -2908 1635
rect -2874 1601 -2858 1635
rect -2806 1601 -2790 1635
rect -2756 1601 -2740 1635
rect -2688 1601 -2672 1635
rect -2638 1601 -2622 1635
rect -2570 1601 -2554 1635
rect -2520 1601 -2504 1635
rect -2452 1601 -2436 1635
rect -2402 1601 -2386 1635
rect -2334 1601 -2318 1635
rect -2284 1601 -2268 1635
rect -2216 1601 -2200 1635
rect -2166 1601 -2150 1635
rect -2098 1601 -2082 1635
rect -2048 1601 -2032 1635
rect -1980 1601 -1964 1635
rect -1930 1601 -1914 1635
rect -1862 1601 -1846 1635
rect -1812 1601 -1796 1635
rect -1744 1601 -1728 1635
rect -1694 1601 -1678 1635
rect -1626 1601 -1610 1635
rect -1576 1601 -1560 1635
rect -1508 1601 -1492 1635
rect -1458 1601 -1442 1635
rect -1390 1601 -1374 1635
rect -1340 1601 -1324 1635
rect -1272 1601 -1256 1635
rect -1222 1601 -1206 1635
rect -1154 1601 -1138 1635
rect -1104 1601 -1088 1635
rect -1036 1601 -1020 1635
rect -986 1601 -970 1635
rect -918 1601 -902 1635
rect -868 1601 -852 1635
rect -800 1601 -784 1635
rect -750 1601 -734 1635
rect -682 1601 -666 1635
rect -632 1601 -616 1635
rect -564 1601 -548 1635
rect -514 1601 -498 1635
rect -446 1601 -430 1635
rect -396 1601 -380 1635
rect -328 1601 -312 1635
rect -278 1601 -262 1635
rect -210 1601 -194 1635
rect -160 1601 -144 1635
rect -92 1601 -76 1635
rect -42 1601 -26 1635
rect 26 1601 42 1635
rect 76 1601 92 1635
rect 144 1601 160 1635
rect 194 1601 210 1635
rect 262 1601 278 1635
rect 312 1601 328 1635
rect 380 1601 396 1635
rect 430 1601 446 1635
rect 498 1601 514 1635
rect 548 1601 564 1635
rect 616 1601 632 1635
rect 666 1601 682 1635
rect 734 1601 750 1635
rect 784 1601 800 1635
rect 852 1601 868 1635
rect 902 1601 918 1635
rect 970 1601 986 1635
rect 1020 1601 1036 1635
rect 1088 1601 1104 1635
rect 1138 1601 1154 1635
rect 1206 1601 1222 1635
rect 1256 1601 1272 1635
rect 1324 1601 1340 1635
rect 1374 1601 1390 1635
rect 1442 1601 1458 1635
rect 1492 1601 1508 1635
rect 1560 1601 1576 1635
rect 1610 1601 1626 1635
rect 1678 1601 1694 1635
rect 1728 1601 1744 1635
rect 1796 1601 1812 1635
rect 1846 1601 1862 1635
rect 1914 1601 1930 1635
rect 1964 1601 1980 1635
rect 2032 1601 2048 1635
rect 2082 1601 2098 1635
rect 2150 1601 2166 1635
rect 2200 1601 2216 1635
rect 2268 1601 2284 1635
rect 2318 1601 2334 1635
rect 2386 1601 2402 1635
rect 2436 1601 2452 1635
rect 2504 1601 2520 1635
rect 2554 1601 2570 1635
rect 2622 1601 2638 1635
rect 2672 1601 2688 1635
rect 2740 1601 2756 1635
rect 2790 1601 2806 1635
rect 2858 1601 2874 1635
rect 2908 1601 2924 1635
rect -2967 1542 -2933 1558
rect -2967 950 -2933 966
rect -2849 1542 -2815 1558
rect -2849 950 -2815 966
rect -2731 1542 -2697 1558
rect -2731 950 -2697 966
rect -2613 1542 -2579 1558
rect -2613 950 -2579 966
rect -2495 1542 -2461 1558
rect -2495 950 -2461 966
rect -2377 1542 -2343 1558
rect -2377 950 -2343 966
rect -2259 1542 -2225 1558
rect -2259 950 -2225 966
rect -2141 1542 -2107 1558
rect -2141 950 -2107 966
rect -2023 1542 -1989 1558
rect -2023 950 -1989 966
rect -1905 1542 -1871 1558
rect -1905 950 -1871 966
rect -1787 1542 -1753 1558
rect -1787 950 -1753 966
rect -1669 1542 -1635 1558
rect -1669 950 -1635 966
rect -1551 1542 -1517 1558
rect -1551 950 -1517 966
rect -1433 1542 -1399 1558
rect -1433 950 -1399 966
rect -1315 1542 -1281 1558
rect -1315 950 -1281 966
rect -1197 1542 -1163 1558
rect -1197 950 -1163 966
rect -1079 1542 -1045 1558
rect -1079 950 -1045 966
rect -961 1542 -927 1558
rect -961 950 -927 966
rect -843 1542 -809 1558
rect -843 950 -809 966
rect -725 1542 -691 1558
rect -725 950 -691 966
rect -607 1542 -573 1558
rect -607 950 -573 966
rect -489 1542 -455 1558
rect -489 950 -455 966
rect -371 1542 -337 1558
rect -371 950 -337 966
rect -253 1542 -219 1558
rect -253 950 -219 966
rect -135 1542 -101 1558
rect -135 950 -101 966
rect -17 1542 17 1558
rect -17 950 17 966
rect 101 1542 135 1558
rect 101 950 135 966
rect 219 1542 253 1558
rect 219 950 253 966
rect 337 1542 371 1558
rect 337 950 371 966
rect 455 1542 489 1558
rect 455 950 489 966
rect 573 1542 607 1558
rect 573 950 607 966
rect 691 1542 725 1558
rect 691 950 725 966
rect 809 1542 843 1558
rect 809 950 843 966
rect 927 1542 961 1558
rect 927 950 961 966
rect 1045 1542 1079 1558
rect 1045 950 1079 966
rect 1163 1542 1197 1558
rect 1163 950 1197 966
rect 1281 1542 1315 1558
rect 1281 950 1315 966
rect 1399 1542 1433 1558
rect 1399 950 1433 966
rect 1517 1542 1551 1558
rect 1517 950 1551 966
rect 1635 1542 1669 1558
rect 1635 950 1669 966
rect 1753 1542 1787 1558
rect 1753 950 1787 966
rect 1871 1542 1905 1558
rect 1871 950 1905 966
rect 1989 1542 2023 1558
rect 1989 950 2023 966
rect 2107 1542 2141 1558
rect 2107 950 2141 966
rect 2225 1542 2259 1558
rect 2225 950 2259 966
rect 2343 1542 2377 1558
rect 2343 950 2377 966
rect 2461 1542 2495 1558
rect 2461 950 2495 966
rect 2579 1542 2613 1558
rect 2579 950 2613 966
rect 2697 1542 2731 1558
rect 2697 950 2731 966
rect 2815 1542 2849 1558
rect 2815 950 2849 966
rect 2933 1542 2967 1558
rect 2933 950 2967 966
rect -2924 873 -2908 907
rect -2874 873 -2858 907
rect -2806 873 -2790 907
rect -2756 873 -2740 907
rect -2688 873 -2672 907
rect -2638 873 -2622 907
rect -2570 873 -2554 907
rect -2520 873 -2504 907
rect -2452 873 -2436 907
rect -2402 873 -2386 907
rect -2334 873 -2318 907
rect -2284 873 -2268 907
rect -2216 873 -2200 907
rect -2166 873 -2150 907
rect -2098 873 -2082 907
rect -2048 873 -2032 907
rect -1980 873 -1964 907
rect -1930 873 -1914 907
rect -1862 873 -1846 907
rect -1812 873 -1796 907
rect -1744 873 -1728 907
rect -1694 873 -1678 907
rect -1626 873 -1610 907
rect -1576 873 -1560 907
rect -1508 873 -1492 907
rect -1458 873 -1442 907
rect -1390 873 -1374 907
rect -1340 873 -1324 907
rect -1272 873 -1256 907
rect -1222 873 -1206 907
rect -1154 873 -1138 907
rect -1104 873 -1088 907
rect -1036 873 -1020 907
rect -986 873 -970 907
rect -918 873 -902 907
rect -868 873 -852 907
rect -800 873 -784 907
rect -750 873 -734 907
rect -682 873 -666 907
rect -632 873 -616 907
rect -564 873 -548 907
rect -514 873 -498 907
rect -446 873 -430 907
rect -396 873 -380 907
rect -328 873 -312 907
rect -278 873 -262 907
rect -210 873 -194 907
rect -160 873 -144 907
rect -92 873 -76 907
rect -42 873 -26 907
rect 26 873 42 907
rect 76 873 92 907
rect 144 873 160 907
rect 194 873 210 907
rect 262 873 278 907
rect 312 873 328 907
rect 380 873 396 907
rect 430 873 446 907
rect 498 873 514 907
rect 548 873 564 907
rect 616 873 632 907
rect 666 873 682 907
rect 734 873 750 907
rect 784 873 800 907
rect 852 873 868 907
rect 902 873 918 907
rect 970 873 986 907
rect 1020 873 1036 907
rect 1088 873 1104 907
rect 1138 873 1154 907
rect 1206 873 1222 907
rect 1256 873 1272 907
rect 1324 873 1340 907
rect 1374 873 1390 907
rect 1442 873 1458 907
rect 1492 873 1508 907
rect 1560 873 1576 907
rect 1610 873 1626 907
rect 1678 873 1694 907
rect 1728 873 1744 907
rect 1796 873 1812 907
rect 1846 873 1862 907
rect 1914 873 1930 907
rect 1964 873 1980 907
rect 2032 873 2048 907
rect 2082 873 2098 907
rect 2150 873 2166 907
rect 2200 873 2216 907
rect 2268 873 2284 907
rect 2318 873 2334 907
rect 2386 873 2402 907
rect 2436 873 2452 907
rect 2504 873 2520 907
rect 2554 873 2570 907
rect 2622 873 2638 907
rect 2672 873 2688 907
rect 2740 873 2756 907
rect 2790 873 2806 907
rect 2858 873 2874 907
rect 2908 873 2924 907
rect -2924 765 -2908 799
rect -2874 765 -2858 799
rect -2806 765 -2790 799
rect -2756 765 -2740 799
rect -2688 765 -2672 799
rect -2638 765 -2622 799
rect -2570 765 -2554 799
rect -2520 765 -2504 799
rect -2452 765 -2436 799
rect -2402 765 -2386 799
rect -2334 765 -2318 799
rect -2284 765 -2268 799
rect -2216 765 -2200 799
rect -2166 765 -2150 799
rect -2098 765 -2082 799
rect -2048 765 -2032 799
rect -1980 765 -1964 799
rect -1930 765 -1914 799
rect -1862 765 -1846 799
rect -1812 765 -1796 799
rect -1744 765 -1728 799
rect -1694 765 -1678 799
rect -1626 765 -1610 799
rect -1576 765 -1560 799
rect -1508 765 -1492 799
rect -1458 765 -1442 799
rect -1390 765 -1374 799
rect -1340 765 -1324 799
rect -1272 765 -1256 799
rect -1222 765 -1206 799
rect -1154 765 -1138 799
rect -1104 765 -1088 799
rect -1036 765 -1020 799
rect -986 765 -970 799
rect -918 765 -902 799
rect -868 765 -852 799
rect -800 765 -784 799
rect -750 765 -734 799
rect -682 765 -666 799
rect -632 765 -616 799
rect -564 765 -548 799
rect -514 765 -498 799
rect -446 765 -430 799
rect -396 765 -380 799
rect -328 765 -312 799
rect -278 765 -262 799
rect -210 765 -194 799
rect -160 765 -144 799
rect -92 765 -76 799
rect -42 765 -26 799
rect 26 765 42 799
rect 76 765 92 799
rect 144 765 160 799
rect 194 765 210 799
rect 262 765 278 799
rect 312 765 328 799
rect 380 765 396 799
rect 430 765 446 799
rect 498 765 514 799
rect 548 765 564 799
rect 616 765 632 799
rect 666 765 682 799
rect 734 765 750 799
rect 784 765 800 799
rect 852 765 868 799
rect 902 765 918 799
rect 970 765 986 799
rect 1020 765 1036 799
rect 1088 765 1104 799
rect 1138 765 1154 799
rect 1206 765 1222 799
rect 1256 765 1272 799
rect 1324 765 1340 799
rect 1374 765 1390 799
rect 1442 765 1458 799
rect 1492 765 1508 799
rect 1560 765 1576 799
rect 1610 765 1626 799
rect 1678 765 1694 799
rect 1728 765 1744 799
rect 1796 765 1812 799
rect 1846 765 1862 799
rect 1914 765 1930 799
rect 1964 765 1980 799
rect 2032 765 2048 799
rect 2082 765 2098 799
rect 2150 765 2166 799
rect 2200 765 2216 799
rect 2268 765 2284 799
rect 2318 765 2334 799
rect 2386 765 2402 799
rect 2436 765 2452 799
rect 2504 765 2520 799
rect 2554 765 2570 799
rect 2622 765 2638 799
rect 2672 765 2688 799
rect 2740 765 2756 799
rect 2790 765 2806 799
rect 2858 765 2874 799
rect 2908 765 2924 799
rect -2967 706 -2933 722
rect -2967 114 -2933 130
rect -2849 706 -2815 722
rect -2849 114 -2815 130
rect -2731 706 -2697 722
rect -2731 114 -2697 130
rect -2613 706 -2579 722
rect -2613 114 -2579 130
rect -2495 706 -2461 722
rect -2495 114 -2461 130
rect -2377 706 -2343 722
rect -2377 114 -2343 130
rect -2259 706 -2225 722
rect -2259 114 -2225 130
rect -2141 706 -2107 722
rect -2141 114 -2107 130
rect -2023 706 -1989 722
rect -2023 114 -1989 130
rect -1905 706 -1871 722
rect -1905 114 -1871 130
rect -1787 706 -1753 722
rect -1787 114 -1753 130
rect -1669 706 -1635 722
rect -1669 114 -1635 130
rect -1551 706 -1517 722
rect -1551 114 -1517 130
rect -1433 706 -1399 722
rect -1433 114 -1399 130
rect -1315 706 -1281 722
rect -1315 114 -1281 130
rect -1197 706 -1163 722
rect -1197 114 -1163 130
rect -1079 706 -1045 722
rect -1079 114 -1045 130
rect -961 706 -927 722
rect -961 114 -927 130
rect -843 706 -809 722
rect -843 114 -809 130
rect -725 706 -691 722
rect -725 114 -691 130
rect -607 706 -573 722
rect -607 114 -573 130
rect -489 706 -455 722
rect -489 114 -455 130
rect -371 706 -337 722
rect -371 114 -337 130
rect -253 706 -219 722
rect -253 114 -219 130
rect -135 706 -101 722
rect -135 114 -101 130
rect -17 706 17 722
rect -17 114 17 130
rect 101 706 135 722
rect 101 114 135 130
rect 219 706 253 722
rect 219 114 253 130
rect 337 706 371 722
rect 337 114 371 130
rect 455 706 489 722
rect 455 114 489 130
rect 573 706 607 722
rect 573 114 607 130
rect 691 706 725 722
rect 691 114 725 130
rect 809 706 843 722
rect 809 114 843 130
rect 927 706 961 722
rect 927 114 961 130
rect 1045 706 1079 722
rect 1045 114 1079 130
rect 1163 706 1197 722
rect 1163 114 1197 130
rect 1281 706 1315 722
rect 1281 114 1315 130
rect 1399 706 1433 722
rect 1399 114 1433 130
rect 1517 706 1551 722
rect 1517 114 1551 130
rect 1635 706 1669 722
rect 1635 114 1669 130
rect 1753 706 1787 722
rect 1753 114 1787 130
rect 1871 706 1905 722
rect 1871 114 1905 130
rect 1989 706 2023 722
rect 1989 114 2023 130
rect 2107 706 2141 722
rect 2107 114 2141 130
rect 2225 706 2259 722
rect 2225 114 2259 130
rect 2343 706 2377 722
rect 2343 114 2377 130
rect 2461 706 2495 722
rect 2461 114 2495 130
rect 2579 706 2613 722
rect 2579 114 2613 130
rect 2697 706 2731 722
rect 2697 114 2731 130
rect 2815 706 2849 722
rect 2815 114 2849 130
rect 2933 706 2967 722
rect 2933 114 2967 130
rect -2924 37 -2908 71
rect -2874 37 -2858 71
rect -2806 37 -2790 71
rect -2756 37 -2740 71
rect -2688 37 -2672 71
rect -2638 37 -2622 71
rect -2570 37 -2554 71
rect -2520 37 -2504 71
rect -2452 37 -2436 71
rect -2402 37 -2386 71
rect -2334 37 -2318 71
rect -2284 37 -2268 71
rect -2216 37 -2200 71
rect -2166 37 -2150 71
rect -2098 37 -2082 71
rect -2048 37 -2032 71
rect -1980 37 -1964 71
rect -1930 37 -1914 71
rect -1862 37 -1846 71
rect -1812 37 -1796 71
rect -1744 37 -1728 71
rect -1694 37 -1678 71
rect -1626 37 -1610 71
rect -1576 37 -1560 71
rect -1508 37 -1492 71
rect -1458 37 -1442 71
rect -1390 37 -1374 71
rect -1340 37 -1324 71
rect -1272 37 -1256 71
rect -1222 37 -1206 71
rect -1154 37 -1138 71
rect -1104 37 -1088 71
rect -1036 37 -1020 71
rect -986 37 -970 71
rect -918 37 -902 71
rect -868 37 -852 71
rect -800 37 -784 71
rect -750 37 -734 71
rect -682 37 -666 71
rect -632 37 -616 71
rect -564 37 -548 71
rect -514 37 -498 71
rect -446 37 -430 71
rect -396 37 -380 71
rect -328 37 -312 71
rect -278 37 -262 71
rect -210 37 -194 71
rect -160 37 -144 71
rect -92 37 -76 71
rect -42 37 -26 71
rect 26 37 42 71
rect 76 37 92 71
rect 144 37 160 71
rect 194 37 210 71
rect 262 37 278 71
rect 312 37 328 71
rect 380 37 396 71
rect 430 37 446 71
rect 498 37 514 71
rect 548 37 564 71
rect 616 37 632 71
rect 666 37 682 71
rect 734 37 750 71
rect 784 37 800 71
rect 852 37 868 71
rect 902 37 918 71
rect 970 37 986 71
rect 1020 37 1036 71
rect 1088 37 1104 71
rect 1138 37 1154 71
rect 1206 37 1222 71
rect 1256 37 1272 71
rect 1324 37 1340 71
rect 1374 37 1390 71
rect 1442 37 1458 71
rect 1492 37 1508 71
rect 1560 37 1576 71
rect 1610 37 1626 71
rect 1678 37 1694 71
rect 1728 37 1744 71
rect 1796 37 1812 71
rect 1846 37 1862 71
rect 1914 37 1930 71
rect 1964 37 1980 71
rect 2032 37 2048 71
rect 2082 37 2098 71
rect 2150 37 2166 71
rect 2200 37 2216 71
rect 2268 37 2284 71
rect 2318 37 2334 71
rect 2386 37 2402 71
rect 2436 37 2452 71
rect 2504 37 2520 71
rect 2554 37 2570 71
rect 2622 37 2638 71
rect 2672 37 2688 71
rect 2740 37 2756 71
rect 2790 37 2806 71
rect 2858 37 2874 71
rect 2908 37 2924 71
rect -2924 -71 -2908 -37
rect -2874 -71 -2858 -37
rect -2806 -71 -2790 -37
rect -2756 -71 -2740 -37
rect -2688 -71 -2672 -37
rect -2638 -71 -2622 -37
rect -2570 -71 -2554 -37
rect -2520 -71 -2504 -37
rect -2452 -71 -2436 -37
rect -2402 -71 -2386 -37
rect -2334 -71 -2318 -37
rect -2284 -71 -2268 -37
rect -2216 -71 -2200 -37
rect -2166 -71 -2150 -37
rect -2098 -71 -2082 -37
rect -2048 -71 -2032 -37
rect -1980 -71 -1964 -37
rect -1930 -71 -1914 -37
rect -1862 -71 -1846 -37
rect -1812 -71 -1796 -37
rect -1744 -71 -1728 -37
rect -1694 -71 -1678 -37
rect -1626 -71 -1610 -37
rect -1576 -71 -1560 -37
rect -1508 -71 -1492 -37
rect -1458 -71 -1442 -37
rect -1390 -71 -1374 -37
rect -1340 -71 -1324 -37
rect -1272 -71 -1256 -37
rect -1222 -71 -1206 -37
rect -1154 -71 -1138 -37
rect -1104 -71 -1088 -37
rect -1036 -71 -1020 -37
rect -986 -71 -970 -37
rect -918 -71 -902 -37
rect -868 -71 -852 -37
rect -800 -71 -784 -37
rect -750 -71 -734 -37
rect -682 -71 -666 -37
rect -632 -71 -616 -37
rect -564 -71 -548 -37
rect -514 -71 -498 -37
rect -446 -71 -430 -37
rect -396 -71 -380 -37
rect -328 -71 -312 -37
rect -278 -71 -262 -37
rect -210 -71 -194 -37
rect -160 -71 -144 -37
rect -92 -71 -76 -37
rect -42 -71 -26 -37
rect 26 -71 42 -37
rect 76 -71 92 -37
rect 144 -71 160 -37
rect 194 -71 210 -37
rect 262 -71 278 -37
rect 312 -71 328 -37
rect 380 -71 396 -37
rect 430 -71 446 -37
rect 498 -71 514 -37
rect 548 -71 564 -37
rect 616 -71 632 -37
rect 666 -71 682 -37
rect 734 -71 750 -37
rect 784 -71 800 -37
rect 852 -71 868 -37
rect 902 -71 918 -37
rect 970 -71 986 -37
rect 1020 -71 1036 -37
rect 1088 -71 1104 -37
rect 1138 -71 1154 -37
rect 1206 -71 1222 -37
rect 1256 -71 1272 -37
rect 1324 -71 1340 -37
rect 1374 -71 1390 -37
rect 1442 -71 1458 -37
rect 1492 -71 1508 -37
rect 1560 -71 1576 -37
rect 1610 -71 1626 -37
rect 1678 -71 1694 -37
rect 1728 -71 1744 -37
rect 1796 -71 1812 -37
rect 1846 -71 1862 -37
rect 1914 -71 1930 -37
rect 1964 -71 1980 -37
rect 2032 -71 2048 -37
rect 2082 -71 2098 -37
rect 2150 -71 2166 -37
rect 2200 -71 2216 -37
rect 2268 -71 2284 -37
rect 2318 -71 2334 -37
rect 2386 -71 2402 -37
rect 2436 -71 2452 -37
rect 2504 -71 2520 -37
rect 2554 -71 2570 -37
rect 2622 -71 2638 -37
rect 2672 -71 2688 -37
rect 2740 -71 2756 -37
rect 2790 -71 2806 -37
rect 2858 -71 2874 -37
rect 2908 -71 2924 -37
rect -2967 -130 -2933 -114
rect -2967 -722 -2933 -706
rect -2849 -130 -2815 -114
rect -2849 -722 -2815 -706
rect -2731 -130 -2697 -114
rect -2731 -722 -2697 -706
rect -2613 -130 -2579 -114
rect -2613 -722 -2579 -706
rect -2495 -130 -2461 -114
rect -2495 -722 -2461 -706
rect -2377 -130 -2343 -114
rect -2377 -722 -2343 -706
rect -2259 -130 -2225 -114
rect -2259 -722 -2225 -706
rect -2141 -130 -2107 -114
rect -2141 -722 -2107 -706
rect -2023 -130 -1989 -114
rect -2023 -722 -1989 -706
rect -1905 -130 -1871 -114
rect -1905 -722 -1871 -706
rect -1787 -130 -1753 -114
rect -1787 -722 -1753 -706
rect -1669 -130 -1635 -114
rect -1669 -722 -1635 -706
rect -1551 -130 -1517 -114
rect -1551 -722 -1517 -706
rect -1433 -130 -1399 -114
rect -1433 -722 -1399 -706
rect -1315 -130 -1281 -114
rect -1315 -722 -1281 -706
rect -1197 -130 -1163 -114
rect -1197 -722 -1163 -706
rect -1079 -130 -1045 -114
rect -1079 -722 -1045 -706
rect -961 -130 -927 -114
rect -961 -722 -927 -706
rect -843 -130 -809 -114
rect -843 -722 -809 -706
rect -725 -130 -691 -114
rect -725 -722 -691 -706
rect -607 -130 -573 -114
rect -607 -722 -573 -706
rect -489 -130 -455 -114
rect -489 -722 -455 -706
rect -371 -130 -337 -114
rect -371 -722 -337 -706
rect -253 -130 -219 -114
rect -253 -722 -219 -706
rect -135 -130 -101 -114
rect -135 -722 -101 -706
rect -17 -130 17 -114
rect -17 -722 17 -706
rect 101 -130 135 -114
rect 101 -722 135 -706
rect 219 -130 253 -114
rect 219 -722 253 -706
rect 337 -130 371 -114
rect 337 -722 371 -706
rect 455 -130 489 -114
rect 455 -722 489 -706
rect 573 -130 607 -114
rect 573 -722 607 -706
rect 691 -130 725 -114
rect 691 -722 725 -706
rect 809 -130 843 -114
rect 809 -722 843 -706
rect 927 -130 961 -114
rect 927 -722 961 -706
rect 1045 -130 1079 -114
rect 1045 -722 1079 -706
rect 1163 -130 1197 -114
rect 1163 -722 1197 -706
rect 1281 -130 1315 -114
rect 1281 -722 1315 -706
rect 1399 -130 1433 -114
rect 1399 -722 1433 -706
rect 1517 -130 1551 -114
rect 1517 -722 1551 -706
rect 1635 -130 1669 -114
rect 1635 -722 1669 -706
rect 1753 -130 1787 -114
rect 1753 -722 1787 -706
rect 1871 -130 1905 -114
rect 1871 -722 1905 -706
rect 1989 -130 2023 -114
rect 1989 -722 2023 -706
rect 2107 -130 2141 -114
rect 2107 -722 2141 -706
rect 2225 -130 2259 -114
rect 2225 -722 2259 -706
rect 2343 -130 2377 -114
rect 2343 -722 2377 -706
rect 2461 -130 2495 -114
rect 2461 -722 2495 -706
rect 2579 -130 2613 -114
rect 2579 -722 2613 -706
rect 2697 -130 2731 -114
rect 2697 -722 2731 -706
rect 2815 -130 2849 -114
rect 2815 -722 2849 -706
rect 2933 -130 2967 -114
rect 2933 -722 2967 -706
rect -2924 -799 -2908 -765
rect -2874 -799 -2858 -765
rect -2806 -799 -2790 -765
rect -2756 -799 -2740 -765
rect -2688 -799 -2672 -765
rect -2638 -799 -2622 -765
rect -2570 -799 -2554 -765
rect -2520 -799 -2504 -765
rect -2452 -799 -2436 -765
rect -2402 -799 -2386 -765
rect -2334 -799 -2318 -765
rect -2284 -799 -2268 -765
rect -2216 -799 -2200 -765
rect -2166 -799 -2150 -765
rect -2098 -799 -2082 -765
rect -2048 -799 -2032 -765
rect -1980 -799 -1964 -765
rect -1930 -799 -1914 -765
rect -1862 -799 -1846 -765
rect -1812 -799 -1796 -765
rect -1744 -799 -1728 -765
rect -1694 -799 -1678 -765
rect -1626 -799 -1610 -765
rect -1576 -799 -1560 -765
rect -1508 -799 -1492 -765
rect -1458 -799 -1442 -765
rect -1390 -799 -1374 -765
rect -1340 -799 -1324 -765
rect -1272 -799 -1256 -765
rect -1222 -799 -1206 -765
rect -1154 -799 -1138 -765
rect -1104 -799 -1088 -765
rect -1036 -799 -1020 -765
rect -986 -799 -970 -765
rect -918 -799 -902 -765
rect -868 -799 -852 -765
rect -800 -799 -784 -765
rect -750 -799 -734 -765
rect -682 -799 -666 -765
rect -632 -799 -616 -765
rect -564 -799 -548 -765
rect -514 -799 -498 -765
rect -446 -799 -430 -765
rect -396 -799 -380 -765
rect -328 -799 -312 -765
rect -278 -799 -262 -765
rect -210 -799 -194 -765
rect -160 -799 -144 -765
rect -92 -799 -76 -765
rect -42 -799 -26 -765
rect 26 -799 42 -765
rect 76 -799 92 -765
rect 144 -799 160 -765
rect 194 -799 210 -765
rect 262 -799 278 -765
rect 312 -799 328 -765
rect 380 -799 396 -765
rect 430 -799 446 -765
rect 498 -799 514 -765
rect 548 -799 564 -765
rect 616 -799 632 -765
rect 666 -799 682 -765
rect 734 -799 750 -765
rect 784 -799 800 -765
rect 852 -799 868 -765
rect 902 -799 918 -765
rect 970 -799 986 -765
rect 1020 -799 1036 -765
rect 1088 -799 1104 -765
rect 1138 -799 1154 -765
rect 1206 -799 1222 -765
rect 1256 -799 1272 -765
rect 1324 -799 1340 -765
rect 1374 -799 1390 -765
rect 1442 -799 1458 -765
rect 1492 -799 1508 -765
rect 1560 -799 1576 -765
rect 1610 -799 1626 -765
rect 1678 -799 1694 -765
rect 1728 -799 1744 -765
rect 1796 -799 1812 -765
rect 1846 -799 1862 -765
rect 1914 -799 1930 -765
rect 1964 -799 1980 -765
rect 2032 -799 2048 -765
rect 2082 -799 2098 -765
rect 2150 -799 2166 -765
rect 2200 -799 2216 -765
rect 2268 -799 2284 -765
rect 2318 -799 2334 -765
rect 2386 -799 2402 -765
rect 2436 -799 2452 -765
rect 2504 -799 2520 -765
rect 2554 -799 2570 -765
rect 2622 -799 2638 -765
rect 2672 -799 2688 -765
rect 2740 -799 2756 -765
rect 2790 -799 2806 -765
rect 2858 -799 2874 -765
rect 2908 -799 2924 -765
rect -2924 -907 -2908 -873
rect -2874 -907 -2858 -873
rect -2806 -907 -2790 -873
rect -2756 -907 -2740 -873
rect -2688 -907 -2672 -873
rect -2638 -907 -2622 -873
rect -2570 -907 -2554 -873
rect -2520 -907 -2504 -873
rect -2452 -907 -2436 -873
rect -2402 -907 -2386 -873
rect -2334 -907 -2318 -873
rect -2284 -907 -2268 -873
rect -2216 -907 -2200 -873
rect -2166 -907 -2150 -873
rect -2098 -907 -2082 -873
rect -2048 -907 -2032 -873
rect -1980 -907 -1964 -873
rect -1930 -907 -1914 -873
rect -1862 -907 -1846 -873
rect -1812 -907 -1796 -873
rect -1744 -907 -1728 -873
rect -1694 -907 -1678 -873
rect -1626 -907 -1610 -873
rect -1576 -907 -1560 -873
rect -1508 -907 -1492 -873
rect -1458 -907 -1442 -873
rect -1390 -907 -1374 -873
rect -1340 -907 -1324 -873
rect -1272 -907 -1256 -873
rect -1222 -907 -1206 -873
rect -1154 -907 -1138 -873
rect -1104 -907 -1088 -873
rect -1036 -907 -1020 -873
rect -986 -907 -970 -873
rect -918 -907 -902 -873
rect -868 -907 -852 -873
rect -800 -907 -784 -873
rect -750 -907 -734 -873
rect -682 -907 -666 -873
rect -632 -907 -616 -873
rect -564 -907 -548 -873
rect -514 -907 -498 -873
rect -446 -907 -430 -873
rect -396 -907 -380 -873
rect -328 -907 -312 -873
rect -278 -907 -262 -873
rect -210 -907 -194 -873
rect -160 -907 -144 -873
rect -92 -907 -76 -873
rect -42 -907 -26 -873
rect 26 -907 42 -873
rect 76 -907 92 -873
rect 144 -907 160 -873
rect 194 -907 210 -873
rect 262 -907 278 -873
rect 312 -907 328 -873
rect 380 -907 396 -873
rect 430 -907 446 -873
rect 498 -907 514 -873
rect 548 -907 564 -873
rect 616 -907 632 -873
rect 666 -907 682 -873
rect 734 -907 750 -873
rect 784 -907 800 -873
rect 852 -907 868 -873
rect 902 -907 918 -873
rect 970 -907 986 -873
rect 1020 -907 1036 -873
rect 1088 -907 1104 -873
rect 1138 -907 1154 -873
rect 1206 -907 1222 -873
rect 1256 -907 1272 -873
rect 1324 -907 1340 -873
rect 1374 -907 1390 -873
rect 1442 -907 1458 -873
rect 1492 -907 1508 -873
rect 1560 -907 1576 -873
rect 1610 -907 1626 -873
rect 1678 -907 1694 -873
rect 1728 -907 1744 -873
rect 1796 -907 1812 -873
rect 1846 -907 1862 -873
rect 1914 -907 1930 -873
rect 1964 -907 1980 -873
rect 2032 -907 2048 -873
rect 2082 -907 2098 -873
rect 2150 -907 2166 -873
rect 2200 -907 2216 -873
rect 2268 -907 2284 -873
rect 2318 -907 2334 -873
rect 2386 -907 2402 -873
rect 2436 -907 2452 -873
rect 2504 -907 2520 -873
rect 2554 -907 2570 -873
rect 2622 -907 2638 -873
rect 2672 -907 2688 -873
rect 2740 -907 2756 -873
rect 2790 -907 2806 -873
rect 2858 -907 2874 -873
rect 2908 -907 2924 -873
rect -2967 -966 -2933 -950
rect -2967 -1558 -2933 -1542
rect -2849 -966 -2815 -950
rect -2849 -1558 -2815 -1542
rect -2731 -966 -2697 -950
rect -2731 -1558 -2697 -1542
rect -2613 -966 -2579 -950
rect -2613 -1558 -2579 -1542
rect -2495 -966 -2461 -950
rect -2495 -1558 -2461 -1542
rect -2377 -966 -2343 -950
rect -2377 -1558 -2343 -1542
rect -2259 -966 -2225 -950
rect -2259 -1558 -2225 -1542
rect -2141 -966 -2107 -950
rect -2141 -1558 -2107 -1542
rect -2023 -966 -1989 -950
rect -2023 -1558 -1989 -1542
rect -1905 -966 -1871 -950
rect -1905 -1558 -1871 -1542
rect -1787 -966 -1753 -950
rect -1787 -1558 -1753 -1542
rect -1669 -966 -1635 -950
rect -1669 -1558 -1635 -1542
rect -1551 -966 -1517 -950
rect -1551 -1558 -1517 -1542
rect -1433 -966 -1399 -950
rect -1433 -1558 -1399 -1542
rect -1315 -966 -1281 -950
rect -1315 -1558 -1281 -1542
rect -1197 -966 -1163 -950
rect -1197 -1558 -1163 -1542
rect -1079 -966 -1045 -950
rect -1079 -1558 -1045 -1542
rect -961 -966 -927 -950
rect -961 -1558 -927 -1542
rect -843 -966 -809 -950
rect -843 -1558 -809 -1542
rect -725 -966 -691 -950
rect -725 -1558 -691 -1542
rect -607 -966 -573 -950
rect -607 -1558 -573 -1542
rect -489 -966 -455 -950
rect -489 -1558 -455 -1542
rect -371 -966 -337 -950
rect -371 -1558 -337 -1542
rect -253 -966 -219 -950
rect -253 -1558 -219 -1542
rect -135 -966 -101 -950
rect -135 -1558 -101 -1542
rect -17 -966 17 -950
rect -17 -1558 17 -1542
rect 101 -966 135 -950
rect 101 -1558 135 -1542
rect 219 -966 253 -950
rect 219 -1558 253 -1542
rect 337 -966 371 -950
rect 337 -1558 371 -1542
rect 455 -966 489 -950
rect 455 -1558 489 -1542
rect 573 -966 607 -950
rect 573 -1558 607 -1542
rect 691 -966 725 -950
rect 691 -1558 725 -1542
rect 809 -966 843 -950
rect 809 -1558 843 -1542
rect 927 -966 961 -950
rect 927 -1558 961 -1542
rect 1045 -966 1079 -950
rect 1045 -1558 1079 -1542
rect 1163 -966 1197 -950
rect 1163 -1558 1197 -1542
rect 1281 -966 1315 -950
rect 1281 -1558 1315 -1542
rect 1399 -966 1433 -950
rect 1399 -1558 1433 -1542
rect 1517 -966 1551 -950
rect 1517 -1558 1551 -1542
rect 1635 -966 1669 -950
rect 1635 -1558 1669 -1542
rect 1753 -966 1787 -950
rect 1753 -1558 1787 -1542
rect 1871 -966 1905 -950
rect 1871 -1558 1905 -1542
rect 1989 -966 2023 -950
rect 1989 -1558 2023 -1542
rect 2107 -966 2141 -950
rect 2107 -1558 2141 -1542
rect 2225 -966 2259 -950
rect 2225 -1558 2259 -1542
rect 2343 -966 2377 -950
rect 2343 -1558 2377 -1542
rect 2461 -966 2495 -950
rect 2461 -1558 2495 -1542
rect 2579 -966 2613 -950
rect 2579 -1558 2613 -1542
rect 2697 -966 2731 -950
rect 2697 -1558 2731 -1542
rect 2815 -966 2849 -950
rect 2815 -1558 2849 -1542
rect 2933 -966 2967 -950
rect 2933 -1558 2967 -1542
rect -2924 -1635 -2908 -1601
rect -2874 -1635 -2858 -1601
rect -2806 -1635 -2790 -1601
rect -2756 -1635 -2740 -1601
rect -2688 -1635 -2672 -1601
rect -2638 -1635 -2622 -1601
rect -2570 -1635 -2554 -1601
rect -2520 -1635 -2504 -1601
rect -2452 -1635 -2436 -1601
rect -2402 -1635 -2386 -1601
rect -2334 -1635 -2318 -1601
rect -2284 -1635 -2268 -1601
rect -2216 -1635 -2200 -1601
rect -2166 -1635 -2150 -1601
rect -2098 -1635 -2082 -1601
rect -2048 -1635 -2032 -1601
rect -1980 -1635 -1964 -1601
rect -1930 -1635 -1914 -1601
rect -1862 -1635 -1846 -1601
rect -1812 -1635 -1796 -1601
rect -1744 -1635 -1728 -1601
rect -1694 -1635 -1678 -1601
rect -1626 -1635 -1610 -1601
rect -1576 -1635 -1560 -1601
rect -1508 -1635 -1492 -1601
rect -1458 -1635 -1442 -1601
rect -1390 -1635 -1374 -1601
rect -1340 -1635 -1324 -1601
rect -1272 -1635 -1256 -1601
rect -1222 -1635 -1206 -1601
rect -1154 -1635 -1138 -1601
rect -1104 -1635 -1088 -1601
rect -1036 -1635 -1020 -1601
rect -986 -1635 -970 -1601
rect -918 -1635 -902 -1601
rect -868 -1635 -852 -1601
rect -800 -1635 -784 -1601
rect -750 -1635 -734 -1601
rect -682 -1635 -666 -1601
rect -632 -1635 -616 -1601
rect -564 -1635 -548 -1601
rect -514 -1635 -498 -1601
rect -446 -1635 -430 -1601
rect -396 -1635 -380 -1601
rect -328 -1635 -312 -1601
rect -278 -1635 -262 -1601
rect -210 -1635 -194 -1601
rect -160 -1635 -144 -1601
rect -92 -1635 -76 -1601
rect -42 -1635 -26 -1601
rect 26 -1635 42 -1601
rect 76 -1635 92 -1601
rect 144 -1635 160 -1601
rect 194 -1635 210 -1601
rect 262 -1635 278 -1601
rect 312 -1635 328 -1601
rect 380 -1635 396 -1601
rect 430 -1635 446 -1601
rect 498 -1635 514 -1601
rect 548 -1635 564 -1601
rect 616 -1635 632 -1601
rect 666 -1635 682 -1601
rect 734 -1635 750 -1601
rect 784 -1635 800 -1601
rect 852 -1635 868 -1601
rect 902 -1635 918 -1601
rect 970 -1635 986 -1601
rect 1020 -1635 1036 -1601
rect 1088 -1635 1104 -1601
rect 1138 -1635 1154 -1601
rect 1206 -1635 1222 -1601
rect 1256 -1635 1272 -1601
rect 1324 -1635 1340 -1601
rect 1374 -1635 1390 -1601
rect 1442 -1635 1458 -1601
rect 1492 -1635 1508 -1601
rect 1560 -1635 1576 -1601
rect 1610 -1635 1626 -1601
rect 1678 -1635 1694 -1601
rect 1728 -1635 1744 -1601
rect 1796 -1635 1812 -1601
rect 1846 -1635 1862 -1601
rect 1914 -1635 1930 -1601
rect 1964 -1635 1980 -1601
rect 2032 -1635 2048 -1601
rect 2082 -1635 2098 -1601
rect 2150 -1635 2166 -1601
rect 2200 -1635 2216 -1601
rect 2268 -1635 2284 -1601
rect 2318 -1635 2334 -1601
rect 2386 -1635 2402 -1601
rect 2436 -1635 2452 -1601
rect 2504 -1635 2520 -1601
rect 2554 -1635 2570 -1601
rect 2622 -1635 2638 -1601
rect 2672 -1635 2688 -1601
rect 2740 -1635 2756 -1601
rect 2790 -1635 2806 -1601
rect 2858 -1635 2874 -1601
rect 2908 -1635 2924 -1601
rect -3081 -1703 -3047 -1641
rect 3047 -1703 3081 -1641
rect -3081 -1737 -2985 -1703
rect 2985 -1737 3081 -1703
<< viali >>
rect -2908 1601 -2874 1635
rect -2790 1601 -2756 1635
rect -2672 1601 -2638 1635
rect -2554 1601 -2520 1635
rect -2436 1601 -2402 1635
rect -2318 1601 -2284 1635
rect -2200 1601 -2166 1635
rect -2082 1601 -2048 1635
rect -1964 1601 -1930 1635
rect -1846 1601 -1812 1635
rect -1728 1601 -1694 1635
rect -1610 1601 -1576 1635
rect -1492 1601 -1458 1635
rect -1374 1601 -1340 1635
rect -1256 1601 -1222 1635
rect -1138 1601 -1104 1635
rect -1020 1601 -986 1635
rect -902 1601 -868 1635
rect -784 1601 -750 1635
rect -666 1601 -632 1635
rect -548 1601 -514 1635
rect -430 1601 -396 1635
rect -312 1601 -278 1635
rect -194 1601 -160 1635
rect -76 1601 -42 1635
rect 42 1601 76 1635
rect 160 1601 194 1635
rect 278 1601 312 1635
rect 396 1601 430 1635
rect 514 1601 548 1635
rect 632 1601 666 1635
rect 750 1601 784 1635
rect 868 1601 902 1635
rect 986 1601 1020 1635
rect 1104 1601 1138 1635
rect 1222 1601 1256 1635
rect 1340 1601 1374 1635
rect 1458 1601 1492 1635
rect 1576 1601 1610 1635
rect 1694 1601 1728 1635
rect 1812 1601 1846 1635
rect 1930 1601 1964 1635
rect 2048 1601 2082 1635
rect 2166 1601 2200 1635
rect 2284 1601 2318 1635
rect 2402 1601 2436 1635
rect 2520 1601 2554 1635
rect 2638 1601 2672 1635
rect 2756 1601 2790 1635
rect 2874 1601 2908 1635
rect -2967 966 -2933 1542
rect -2849 966 -2815 1542
rect -2731 966 -2697 1542
rect -2613 966 -2579 1542
rect -2495 966 -2461 1542
rect -2377 966 -2343 1542
rect -2259 966 -2225 1542
rect -2141 966 -2107 1542
rect -2023 966 -1989 1542
rect -1905 966 -1871 1542
rect -1787 966 -1753 1542
rect -1669 966 -1635 1542
rect -1551 966 -1517 1542
rect -1433 966 -1399 1542
rect -1315 966 -1281 1542
rect -1197 966 -1163 1542
rect -1079 966 -1045 1542
rect -961 966 -927 1542
rect -843 966 -809 1542
rect -725 966 -691 1542
rect -607 966 -573 1542
rect -489 966 -455 1542
rect -371 966 -337 1542
rect -253 966 -219 1542
rect -135 966 -101 1542
rect -17 966 17 1542
rect 101 966 135 1542
rect 219 966 253 1542
rect 337 966 371 1542
rect 455 966 489 1542
rect 573 966 607 1542
rect 691 966 725 1542
rect 809 966 843 1542
rect 927 966 961 1542
rect 1045 966 1079 1542
rect 1163 966 1197 1542
rect 1281 966 1315 1542
rect 1399 966 1433 1542
rect 1517 966 1551 1542
rect 1635 966 1669 1542
rect 1753 966 1787 1542
rect 1871 966 1905 1542
rect 1989 966 2023 1542
rect 2107 966 2141 1542
rect 2225 966 2259 1542
rect 2343 966 2377 1542
rect 2461 966 2495 1542
rect 2579 966 2613 1542
rect 2697 966 2731 1542
rect 2815 966 2849 1542
rect 2933 966 2967 1542
rect -2908 873 -2874 907
rect -2790 873 -2756 907
rect -2672 873 -2638 907
rect -2554 873 -2520 907
rect -2436 873 -2402 907
rect -2318 873 -2284 907
rect -2200 873 -2166 907
rect -2082 873 -2048 907
rect -1964 873 -1930 907
rect -1846 873 -1812 907
rect -1728 873 -1694 907
rect -1610 873 -1576 907
rect -1492 873 -1458 907
rect -1374 873 -1340 907
rect -1256 873 -1222 907
rect -1138 873 -1104 907
rect -1020 873 -986 907
rect -902 873 -868 907
rect -784 873 -750 907
rect -666 873 -632 907
rect -548 873 -514 907
rect -430 873 -396 907
rect -312 873 -278 907
rect -194 873 -160 907
rect -76 873 -42 907
rect 42 873 76 907
rect 160 873 194 907
rect 278 873 312 907
rect 396 873 430 907
rect 514 873 548 907
rect 632 873 666 907
rect 750 873 784 907
rect 868 873 902 907
rect 986 873 1020 907
rect 1104 873 1138 907
rect 1222 873 1256 907
rect 1340 873 1374 907
rect 1458 873 1492 907
rect 1576 873 1610 907
rect 1694 873 1728 907
rect 1812 873 1846 907
rect 1930 873 1964 907
rect 2048 873 2082 907
rect 2166 873 2200 907
rect 2284 873 2318 907
rect 2402 873 2436 907
rect 2520 873 2554 907
rect 2638 873 2672 907
rect 2756 873 2790 907
rect 2874 873 2908 907
rect -2908 765 -2874 799
rect -2790 765 -2756 799
rect -2672 765 -2638 799
rect -2554 765 -2520 799
rect -2436 765 -2402 799
rect -2318 765 -2284 799
rect -2200 765 -2166 799
rect -2082 765 -2048 799
rect -1964 765 -1930 799
rect -1846 765 -1812 799
rect -1728 765 -1694 799
rect -1610 765 -1576 799
rect -1492 765 -1458 799
rect -1374 765 -1340 799
rect -1256 765 -1222 799
rect -1138 765 -1104 799
rect -1020 765 -986 799
rect -902 765 -868 799
rect -784 765 -750 799
rect -666 765 -632 799
rect -548 765 -514 799
rect -430 765 -396 799
rect -312 765 -278 799
rect -194 765 -160 799
rect -76 765 -42 799
rect 42 765 76 799
rect 160 765 194 799
rect 278 765 312 799
rect 396 765 430 799
rect 514 765 548 799
rect 632 765 666 799
rect 750 765 784 799
rect 868 765 902 799
rect 986 765 1020 799
rect 1104 765 1138 799
rect 1222 765 1256 799
rect 1340 765 1374 799
rect 1458 765 1492 799
rect 1576 765 1610 799
rect 1694 765 1728 799
rect 1812 765 1846 799
rect 1930 765 1964 799
rect 2048 765 2082 799
rect 2166 765 2200 799
rect 2284 765 2318 799
rect 2402 765 2436 799
rect 2520 765 2554 799
rect 2638 765 2672 799
rect 2756 765 2790 799
rect 2874 765 2908 799
rect -2967 130 -2933 706
rect -2849 130 -2815 706
rect -2731 130 -2697 706
rect -2613 130 -2579 706
rect -2495 130 -2461 706
rect -2377 130 -2343 706
rect -2259 130 -2225 706
rect -2141 130 -2107 706
rect -2023 130 -1989 706
rect -1905 130 -1871 706
rect -1787 130 -1753 706
rect -1669 130 -1635 706
rect -1551 130 -1517 706
rect -1433 130 -1399 706
rect -1315 130 -1281 706
rect -1197 130 -1163 706
rect -1079 130 -1045 706
rect -961 130 -927 706
rect -843 130 -809 706
rect -725 130 -691 706
rect -607 130 -573 706
rect -489 130 -455 706
rect -371 130 -337 706
rect -253 130 -219 706
rect -135 130 -101 706
rect -17 130 17 706
rect 101 130 135 706
rect 219 130 253 706
rect 337 130 371 706
rect 455 130 489 706
rect 573 130 607 706
rect 691 130 725 706
rect 809 130 843 706
rect 927 130 961 706
rect 1045 130 1079 706
rect 1163 130 1197 706
rect 1281 130 1315 706
rect 1399 130 1433 706
rect 1517 130 1551 706
rect 1635 130 1669 706
rect 1753 130 1787 706
rect 1871 130 1905 706
rect 1989 130 2023 706
rect 2107 130 2141 706
rect 2225 130 2259 706
rect 2343 130 2377 706
rect 2461 130 2495 706
rect 2579 130 2613 706
rect 2697 130 2731 706
rect 2815 130 2849 706
rect 2933 130 2967 706
rect -2908 37 -2874 71
rect -2790 37 -2756 71
rect -2672 37 -2638 71
rect -2554 37 -2520 71
rect -2436 37 -2402 71
rect -2318 37 -2284 71
rect -2200 37 -2166 71
rect -2082 37 -2048 71
rect -1964 37 -1930 71
rect -1846 37 -1812 71
rect -1728 37 -1694 71
rect -1610 37 -1576 71
rect -1492 37 -1458 71
rect -1374 37 -1340 71
rect -1256 37 -1222 71
rect -1138 37 -1104 71
rect -1020 37 -986 71
rect -902 37 -868 71
rect -784 37 -750 71
rect -666 37 -632 71
rect -548 37 -514 71
rect -430 37 -396 71
rect -312 37 -278 71
rect -194 37 -160 71
rect -76 37 -42 71
rect 42 37 76 71
rect 160 37 194 71
rect 278 37 312 71
rect 396 37 430 71
rect 514 37 548 71
rect 632 37 666 71
rect 750 37 784 71
rect 868 37 902 71
rect 986 37 1020 71
rect 1104 37 1138 71
rect 1222 37 1256 71
rect 1340 37 1374 71
rect 1458 37 1492 71
rect 1576 37 1610 71
rect 1694 37 1728 71
rect 1812 37 1846 71
rect 1930 37 1964 71
rect 2048 37 2082 71
rect 2166 37 2200 71
rect 2284 37 2318 71
rect 2402 37 2436 71
rect 2520 37 2554 71
rect 2638 37 2672 71
rect 2756 37 2790 71
rect 2874 37 2908 71
rect -2908 -71 -2874 -37
rect -2790 -71 -2756 -37
rect -2672 -71 -2638 -37
rect -2554 -71 -2520 -37
rect -2436 -71 -2402 -37
rect -2318 -71 -2284 -37
rect -2200 -71 -2166 -37
rect -2082 -71 -2048 -37
rect -1964 -71 -1930 -37
rect -1846 -71 -1812 -37
rect -1728 -71 -1694 -37
rect -1610 -71 -1576 -37
rect -1492 -71 -1458 -37
rect -1374 -71 -1340 -37
rect -1256 -71 -1222 -37
rect -1138 -71 -1104 -37
rect -1020 -71 -986 -37
rect -902 -71 -868 -37
rect -784 -71 -750 -37
rect -666 -71 -632 -37
rect -548 -71 -514 -37
rect -430 -71 -396 -37
rect -312 -71 -278 -37
rect -194 -71 -160 -37
rect -76 -71 -42 -37
rect 42 -71 76 -37
rect 160 -71 194 -37
rect 278 -71 312 -37
rect 396 -71 430 -37
rect 514 -71 548 -37
rect 632 -71 666 -37
rect 750 -71 784 -37
rect 868 -71 902 -37
rect 986 -71 1020 -37
rect 1104 -71 1138 -37
rect 1222 -71 1256 -37
rect 1340 -71 1374 -37
rect 1458 -71 1492 -37
rect 1576 -71 1610 -37
rect 1694 -71 1728 -37
rect 1812 -71 1846 -37
rect 1930 -71 1964 -37
rect 2048 -71 2082 -37
rect 2166 -71 2200 -37
rect 2284 -71 2318 -37
rect 2402 -71 2436 -37
rect 2520 -71 2554 -37
rect 2638 -71 2672 -37
rect 2756 -71 2790 -37
rect 2874 -71 2908 -37
rect -2967 -706 -2933 -130
rect -2849 -706 -2815 -130
rect -2731 -706 -2697 -130
rect -2613 -706 -2579 -130
rect -2495 -706 -2461 -130
rect -2377 -706 -2343 -130
rect -2259 -706 -2225 -130
rect -2141 -706 -2107 -130
rect -2023 -706 -1989 -130
rect -1905 -706 -1871 -130
rect -1787 -706 -1753 -130
rect -1669 -706 -1635 -130
rect -1551 -706 -1517 -130
rect -1433 -706 -1399 -130
rect -1315 -706 -1281 -130
rect -1197 -706 -1163 -130
rect -1079 -706 -1045 -130
rect -961 -706 -927 -130
rect -843 -706 -809 -130
rect -725 -706 -691 -130
rect -607 -706 -573 -130
rect -489 -706 -455 -130
rect -371 -706 -337 -130
rect -253 -706 -219 -130
rect -135 -706 -101 -130
rect -17 -706 17 -130
rect 101 -706 135 -130
rect 219 -706 253 -130
rect 337 -706 371 -130
rect 455 -706 489 -130
rect 573 -706 607 -130
rect 691 -706 725 -130
rect 809 -706 843 -130
rect 927 -706 961 -130
rect 1045 -706 1079 -130
rect 1163 -706 1197 -130
rect 1281 -706 1315 -130
rect 1399 -706 1433 -130
rect 1517 -706 1551 -130
rect 1635 -706 1669 -130
rect 1753 -706 1787 -130
rect 1871 -706 1905 -130
rect 1989 -706 2023 -130
rect 2107 -706 2141 -130
rect 2225 -706 2259 -130
rect 2343 -706 2377 -130
rect 2461 -706 2495 -130
rect 2579 -706 2613 -130
rect 2697 -706 2731 -130
rect 2815 -706 2849 -130
rect 2933 -706 2967 -130
rect -2908 -799 -2874 -765
rect -2790 -799 -2756 -765
rect -2672 -799 -2638 -765
rect -2554 -799 -2520 -765
rect -2436 -799 -2402 -765
rect -2318 -799 -2284 -765
rect -2200 -799 -2166 -765
rect -2082 -799 -2048 -765
rect -1964 -799 -1930 -765
rect -1846 -799 -1812 -765
rect -1728 -799 -1694 -765
rect -1610 -799 -1576 -765
rect -1492 -799 -1458 -765
rect -1374 -799 -1340 -765
rect -1256 -799 -1222 -765
rect -1138 -799 -1104 -765
rect -1020 -799 -986 -765
rect -902 -799 -868 -765
rect -784 -799 -750 -765
rect -666 -799 -632 -765
rect -548 -799 -514 -765
rect -430 -799 -396 -765
rect -312 -799 -278 -765
rect -194 -799 -160 -765
rect -76 -799 -42 -765
rect 42 -799 76 -765
rect 160 -799 194 -765
rect 278 -799 312 -765
rect 396 -799 430 -765
rect 514 -799 548 -765
rect 632 -799 666 -765
rect 750 -799 784 -765
rect 868 -799 902 -765
rect 986 -799 1020 -765
rect 1104 -799 1138 -765
rect 1222 -799 1256 -765
rect 1340 -799 1374 -765
rect 1458 -799 1492 -765
rect 1576 -799 1610 -765
rect 1694 -799 1728 -765
rect 1812 -799 1846 -765
rect 1930 -799 1964 -765
rect 2048 -799 2082 -765
rect 2166 -799 2200 -765
rect 2284 -799 2318 -765
rect 2402 -799 2436 -765
rect 2520 -799 2554 -765
rect 2638 -799 2672 -765
rect 2756 -799 2790 -765
rect 2874 -799 2908 -765
rect -2908 -907 -2874 -873
rect -2790 -907 -2756 -873
rect -2672 -907 -2638 -873
rect -2554 -907 -2520 -873
rect -2436 -907 -2402 -873
rect -2318 -907 -2284 -873
rect -2200 -907 -2166 -873
rect -2082 -907 -2048 -873
rect -1964 -907 -1930 -873
rect -1846 -907 -1812 -873
rect -1728 -907 -1694 -873
rect -1610 -907 -1576 -873
rect -1492 -907 -1458 -873
rect -1374 -907 -1340 -873
rect -1256 -907 -1222 -873
rect -1138 -907 -1104 -873
rect -1020 -907 -986 -873
rect -902 -907 -868 -873
rect -784 -907 -750 -873
rect -666 -907 -632 -873
rect -548 -907 -514 -873
rect -430 -907 -396 -873
rect -312 -907 -278 -873
rect -194 -907 -160 -873
rect -76 -907 -42 -873
rect 42 -907 76 -873
rect 160 -907 194 -873
rect 278 -907 312 -873
rect 396 -907 430 -873
rect 514 -907 548 -873
rect 632 -907 666 -873
rect 750 -907 784 -873
rect 868 -907 902 -873
rect 986 -907 1020 -873
rect 1104 -907 1138 -873
rect 1222 -907 1256 -873
rect 1340 -907 1374 -873
rect 1458 -907 1492 -873
rect 1576 -907 1610 -873
rect 1694 -907 1728 -873
rect 1812 -907 1846 -873
rect 1930 -907 1964 -873
rect 2048 -907 2082 -873
rect 2166 -907 2200 -873
rect 2284 -907 2318 -873
rect 2402 -907 2436 -873
rect 2520 -907 2554 -873
rect 2638 -907 2672 -873
rect 2756 -907 2790 -873
rect 2874 -907 2908 -873
rect -2967 -1542 -2933 -966
rect -2849 -1542 -2815 -966
rect -2731 -1542 -2697 -966
rect -2613 -1542 -2579 -966
rect -2495 -1542 -2461 -966
rect -2377 -1542 -2343 -966
rect -2259 -1542 -2225 -966
rect -2141 -1542 -2107 -966
rect -2023 -1542 -1989 -966
rect -1905 -1542 -1871 -966
rect -1787 -1542 -1753 -966
rect -1669 -1542 -1635 -966
rect -1551 -1542 -1517 -966
rect -1433 -1542 -1399 -966
rect -1315 -1542 -1281 -966
rect -1197 -1542 -1163 -966
rect -1079 -1542 -1045 -966
rect -961 -1542 -927 -966
rect -843 -1542 -809 -966
rect -725 -1542 -691 -966
rect -607 -1542 -573 -966
rect -489 -1542 -455 -966
rect -371 -1542 -337 -966
rect -253 -1542 -219 -966
rect -135 -1542 -101 -966
rect -17 -1542 17 -966
rect 101 -1542 135 -966
rect 219 -1542 253 -966
rect 337 -1542 371 -966
rect 455 -1542 489 -966
rect 573 -1542 607 -966
rect 691 -1542 725 -966
rect 809 -1542 843 -966
rect 927 -1542 961 -966
rect 1045 -1542 1079 -966
rect 1163 -1542 1197 -966
rect 1281 -1542 1315 -966
rect 1399 -1542 1433 -966
rect 1517 -1542 1551 -966
rect 1635 -1542 1669 -966
rect 1753 -1542 1787 -966
rect 1871 -1542 1905 -966
rect 1989 -1542 2023 -966
rect 2107 -1542 2141 -966
rect 2225 -1542 2259 -966
rect 2343 -1542 2377 -966
rect 2461 -1542 2495 -966
rect 2579 -1542 2613 -966
rect 2697 -1542 2731 -966
rect 2815 -1542 2849 -966
rect 2933 -1542 2967 -966
rect -2908 -1635 -2874 -1601
rect -2790 -1635 -2756 -1601
rect -2672 -1635 -2638 -1601
rect -2554 -1635 -2520 -1601
rect -2436 -1635 -2402 -1601
rect -2318 -1635 -2284 -1601
rect -2200 -1635 -2166 -1601
rect -2082 -1635 -2048 -1601
rect -1964 -1635 -1930 -1601
rect -1846 -1635 -1812 -1601
rect -1728 -1635 -1694 -1601
rect -1610 -1635 -1576 -1601
rect -1492 -1635 -1458 -1601
rect -1374 -1635 -1340 -1601
rect -1256 -1635 -1222 -1601
rect -1138 -1635 -1104 -1601
rect -1020 -1635 -986 -1601
rect -902 -1635 -868 -1601
rect -784 -1635 -750 -1601
rect -666 -1635 -632 -1601
rect -548 -1635 -514 -1601
rect -430 -1635 -396 -1601
rect -312 -1635 -278 -1601
rect -194 -1635 -160 -1601
rect -76 -1635 -42 -1601
rect 42 -1635 76 -1601
rect 160 -1635 194 -1601
rect 278 -1635 312 -1601
rect 396 -1635 430 -1601
rect 514 -1635 548 -1601
rect 632 -1635 666 -1601
rect 750 -1635 784 -1601
rect 868 -1635 902 -1601
rect 986 -1635 1020 -1601
rect 1104 -1635 1138 -1601
rect 1222 -1635 1256 -1601
rect 1340 -1635 1374 -1601
rect 1458 -1635 1492 -1601
rect 1576 -1635 1610 -1601
rect 1694 -1635 1728 -1601
rect 1812 -1635 1846 -1601
rect 1930 -1635 1964 -1601
rect 2048 -1635 2082 -1601
rect 2166 -1635 2200 -1601
rect 2284 -1635 2318 -1601
rect 2402 -1635 2436 -1601
rect 2520 -1635 2554 -1601
rect 2638 -1635 2672 -1601
rect 2756 -1635 2790 -1601
rect 2874 -1635 2908 -1601
<< metal1 >>
rect -2920 1635 -2862 1641
rect -2920 1601 -2908 1635
rect -2874 1601 -2862 1635
rect -2920 1595 -2862 1601
rect -2802 1635 -2744 1641
rect -2802 1601 -2790 1635
rect -2756 1601 -2744 1635
rect -2802 1595 -2744 1601
rect -2684 1635 -2626 1641
rect -2684 1601 -2672 1635
rect -2638 1601 -2626 1635
rect -2684 1595 -2626 1601
rect -2566 1635 -2508 1641
rect -2566 1601 -2554 1635
rect -2520 1601 -2508 1635
rect -2566 1595 -2508 1601
rect -2448 1635 -2390 1641
rect -2448 1601 -2436 1635
rect -2402 1601 -2390 1635
rect -2448 1595 -2390 1601
rect -2330 1635 -2272 1641
rect -2330 1601 -2318 1635
rect -2284 1601 -2272 1635
rect -2330 1595 -2272 1601
rect -2212 1635 -2154 1641
rect -2212 1601 -2200 1635
rect -2166 1601 -2154 1635
rect -2212 1595 -2154 1601
rect -2094 1635 -2036 1641
rect -2094 1601 -2082 1635
rect -2048 1601 -2036 1635
rect -2094 1595 -2036 1601
rect -1976 1635 -1918 1641
rect -1976 1601 -1964 1635
rect -1930 1601 -1918 1635
rect -1976 1595 -1918 1601
rect -1858 1635 -1800 1641
rect -1858 1601 -1846 1635
rect -1812 1601 -1800 1635
rect -1858 1595 -1800 1601
rect -1740 1635 -1682 1641
rect -1740 1601 -1728 1635
rect -1694 1601 -1682 1635
rect -1740 1595 -1682 1601
rect -1622 1635 -1564 1641
rect -1622 1601 -1610 1635
rect -1576 1601 -1564 1635
rect -1622 1595 -1564 1601
rect -1504 1635 -1446 1641
rect -1504 1601 -1492 1635
rect -1458 1601 -1446 1635
rect -1504 1595 -1446 1601
rect -1386 1635 -1328 1641
rect -1386 1601 -1374 1635
rect -1340 1601 -1328 1635
rect -1386 1595 -1328 1601
rect -1268 1635 -1210 1641
rect -1268 1601 -1256 1635
rect -1222 1601 -1210 1635
rect -1268 1595 -1210 1601
rect -1150 1635 -1092 1641
rect -1150 1601 -1138 1635
rect -1104 1601 -1092 1635
rect -1150 1595 -1092 1601
rect -1032 1635 -974 1641
rect -1032 1601 -1020 1635
rect -986 1601 -974 1635
rect -1032 1595 -974 1601
rect -914 1635 -856 1641
rect -914 1601 -902 1635
rect -868 1601 -856 1635
rect -914 1595 -856 1601
rect -796 1635 -738 1641
rect -796 1601 -784 1635
rect -750 1601 -738 1635
rect -796 1595 -738 1601
rect -678 1635 -620 1641
rect -678 1601 -666 1635
rect -632 1601 -620 1635
rect -678 1595 -620 1601
rect -560 1635 -502 1641
rect -560 1601 -548 1635
rect -514 1601 -502 1635
rect -560 1595 -502 1601
rect -442 1635 -384 1641
rect -442 1601 -430 1635
rect -396 1601 -384 1635
rect -442 1595 -384 1601
rect -324 1635 -266 1641
rect -324 1601 -312 1635
rect -278 1601 -266 1635
rect -324 1595 -266 1601
rect -206 1635 -148 1641
rect -206 1601 -194 1635
rect -160 1601 -148 1635
rect -206 1595 -148 1601
rect -88 1635 -30 1641
rect -88 1601 -76 1635
rect -42 1601 -30 1635
rect -88 1595 -30 1601
rect 30 1635 88 1641
rect 30 1601 42 1635
rect 76 1601 88 1635
rect 30 1595 88 1601
rect 148 1635 206 1641
rect 148 1601 160 1635
rect 194 1601 206 1635
rect 148 1595 206 1601
rect 266 1635 324 1641
rect 266 1601 278 1635
rect 312 1601 324 1635
rect 266 1595 324 1601
rect 384 1635 442 1641
rect 384 1601 396 1635
rect 430 1601 442 1635
rect 384 1595 442 1601
rect 502 1635 560 1641
rect 502 1601 514 1635
rect 548 1601 560 1635
rect 502 1595 560 1601
rect 620 1635 678 1641
rect 620 1601 632 1635
rect 666 1601 678 1635
rect 620 1595 678 1601
rect 738 1635 796 1641
rect 738 1601 750 1635
rect 784 1601 796 1635
rect 738 1595 796 1601
rect 856 1635 914 1641
rect 856 1601 868 1635
rect 902 1601 914 1635
rect 856 1595 914 1601
rect 974 1635 1032 1641
rect 974 1601 986 1635
rect 1020 1601 1032 1635
rect 974 1595 1032 1601
rect 1092 1635 1150 1641
rect 1092 1601 1104 1635
rect 1138 1601 1150 1635
rect 1092 1595 1150 1601
rect 1210 1635 1268 1641
rect 1210 1601 1222 1635
rect 1256 1601 1268 1635
rect 1210 1595 1268 1601
rect 1328 1635 1386 1641
rect 1328 1601 1340 1635
rect 1374 1601 1386 1635
rect 1328 1595 1386 1601
rect 1446 1635 1504 1641
rect 1446 1601 1458 1635
rect 1492 1601 1504 1635
rect 1446 1595 1504 1601
rect 1564 1635 1622 1641
rect 1564 1601 1576 1635
rect 1610 1601 1622 1635
rect 1564 1595 1622 1601
rect 1682 1635 1740 1641
rect 1682 1601 1694 1635
rect 1728 1601 1740 1635
rect 1682 1595 1740 1601
rect 1800 1635 1858 1641
rect 1800 1601 1812 1635
rect 1846 1601 1858 1635
rect 1800 1595 1858 1601
rect 1918 1635 1976 1641
rect 1918 1601 1930 1635
rect 1964 1601 1976 1635
rect 1918 1595 1976 1601
rect 2036 1635 2094 1641
rect 2036 1601 2048 1635
rect 2082 1601 2094 1635
rect 2036 1595 2094 1601
rect 2154 1635 2212 1641
rect 2154 1601 2166 1635
rect 2200 1601 2212 1635
rect 2154 1595 2212 1601
rect 2272 1635 2330 1641
rect 2272 1601 2284 1635
rect 2318 1601 2330 1635
rect 2272 1595 2330 1601
rect 2390 1635 2448 1641
rect 2390 1601 2402 1635
rect 2436 1601 2448 1635
rect 2390 1595 2448 1601
rect 2508 1635 2566 1641
rect 2508 1601 2520 1635
rect 2554 1601 2566 1635
rect 2508 1595 2566 1601
rect 2626 1635 2684 1641
rect 2626 1601 2638 1635
rect 2672 1601 2684 1635
rect 2626 1595 2684 1601
rect 2744 1635 2802 1641
rect 2744 1601 2756 1635
rect 2790 1601 2802 1635
rect 2744 1595 2802 1601
rect 2862 1635 2920 1641
rect 2862 1601 2874 1635
rect 2908 1601 2920 1635
rect 2862 1595 2920 1601
rect -2973 1542 -2927 1554
rect -2973 966 -2967 1542
rect -2933 966 -2927 1542
rect -2973 954 -2927 966
rect -2855 1542 -2809 1554
rect -2855 966 -2849 1542
rect -2815 966 -2809 1542
rect -2855 954 -2809 966
rect -2737 1542 -2691 1554
rect -2737 966 -2731 1542
rect -2697 966 -2691 1542
rect -2737 954 -2691 966
rect -2619 1542 -2573 1554
rect -2619 966 -2613 1542
rect -2579 966 -2573 1542
rect -2619 954 -2573 966
rect -2501 1542 -2455 1554
rect -2501 966 -2495 1542
rect -2461 966 -2455 1542
rect -2501 954 -2455 966
rect -2383 1542 -2337 1554
rect -2383 966 -2377 1542
rect -2343 966 -2337 1542
rect -2383 954 -2337 966
rect -2265 1542 -2219 1554
rect -2265 966 -2259 1542
rect -2225 966 -2219 1542
rect -2265 954 -2219 966
rect -2147 1542 -2101 1554
rect -2147 966 -2141 1542
rect -2107 966 -2101 1542
rect -2147 954 -2101 966
rect -2029 1542 -1983 1554
rect -2029 966 -2023 1542
rect -1989 966 -1983 1542
rect -2029 954 -1983 966
rect -1911 1542 -1865 1554
rect -1911 966 -1905 1542
rect -1871 966 -1865 1542
rect -1911 954 -1865 966
rect -1793 1542 -1747 1554
rect -1793 966 -1787 1542
rect -1753 966 -1747 1542
rect -1793 954 -1747 966
rect -1675 1542 -1629 1554
rect -1675 966 -1669 1542
rect -1635 966 -1629 1542
rect -1675 954 -1629 966
rect -1557 1542 -1511 1554
rect -1557 966 -1551 1542
rect -1517 966 -1511 1542
rect -1557 954 -1511 966
rect -1439 1542 -1393 1554
rect -1439 966 -1433 1542
rect -1399 966 -1393 1542
rect -1439 954 -1393 966
rect -1321 1542 -1275 1554
rect -1321 966 -1315 1542
rect -1281 966 -1275 1542
rect -1321 954 -1275 966
rect -1203 1542 -1157 1554
rect -1203 966 -1197 1542
rect -1163 966 -1157 1542
rect -1203 954 -1157 966
rect -1085 1542 -1039 1554
rect -1085 966 -1079 1542
rect -1045 966 -1039 1542
rect -1085 954 -1039 966
rect -967 1542 -921 1554
rect -967 966 -961 1542
rect -927 966 -921 1542
rect -967 954 -921 966
rect -849 1542 -803 1554
rect -849 966 -843 1542
rect -809 966 -803 1542
rect -849 954 -803 966
rect -731 1542 -685 1554
rect -731 966 -725 1542
rect -691 966 -685 1542
rect -731 954 -685 966
rect -613 1542 -567 1554
rect -613 966 -607 1542
rect -573 966 -567 1542
rect -613 954 -567 966
rect -495 1542 -449 1554
rect -495 966 -489 1542
rect -455 966 -449 1542
rect -495 954 -449 966
rect -377 1542 -331 1554
rect -377 966 -371 1542
rect -337 966 -331 1542
rect -377 954 -331 966
rect -259 1542 -213 1554
rect -259 966 -253 1542
rect -219 966 -213 1542
rect -259 954 -213 966
rect -141 1542 -95 1554
rect -141 966 -135 1542
rect -101 966 -95 1542
rect -141 954 -95 966
rect -23 1542 23 1554
rect -23 966 -17 1542
rect 17 966 23 1542
rect -23 954 23 966
rect 95 1542 141 1554
rect 95 966 101 1542
rect 135 966 141 1542
rect 95 954 141 966
rect 213 1542 259 1554
rect 213 966 219 1542
rect 253 966 259 1542
rect 213 954 259 966
rect 331 1542 377 1554
rect 331 966 337 1542
rect 371 966 377 1542
rect 331 954 377 966
rect 449 1542 495 1554
rect 449 966 455 1542
rect 489 966 495 1542
rect 449 954 495 966
rect 567 1542 613 1554
rect 567 966 573 1542
rect 607 966 613 1542
rect 567 954 613 966
rect 685 1542 731 1554
rect 685 966 691 1542
rect 725 966 731 1542
rect 685 954 731 966
rect 803 1542 849 1554
rect 803 966 809 1542
rect 843 966 849 1542
rect 803 954 849 966
rect 921 1542 967 1554
rect 921 966 927 1542
rect 961 966 967 1542
rect 921 954 967 966
rect 1039 1542 1085 1554
rect 1039 966 1045 1542
rect 1079 966 1085 1542
rect 1039 954 1085 966
rect 1157 1542 1203 1554
rect 1157 966 1163 1542
rect 1197 966 1203 1542
rect 1157 954 1203 966
rect 1275 1542 1321 1554
rect 1275 966 1281 1542
rect 1315 966 1321 1542
rect 1275 954 1321 966
rect 1393 1542 1439 1554
rect 1393 966 1399 1542
rect 1433 966 1439 1542
rect 1393 954 1439 966
rect 1511 1542 1557 1554
rect 1511 966 1517 1542
rect 1551 966 1557 1542
rect 1511 954 1557 966
rect 1629 1542 1675 1554
rect 1629 966 1635 1542
rect 1669 966 1675 1542
rect 1629 954 1675 966
rect 1747 1542 1793 1554
rect 1747 966 1753 1542
rect 1787 966 1793 1542
rect 1747 954 1793 966
rect 1865 1542 1911 1554
rect 1865 966 1871 1542
rect 1905 966 1911 1542
rect 1865 954 1911 966
rect 1983 1542 2029 1554
rect 1983 966 1989 1542
rect 2023 966 2029 1542
rect 1983 954 2029 966
rect 2101 1542 2147 1554
rect 2101 966 2107 1542
rect 2141 966 2147 1542
rect 2101 954 2147 966
rect 2219 1542 2265 1554
rect 2219 966 2225 1542
rect 2259 966 2265 1542
rect 2219 954 2265 966
rect 2337 1542 2383 1554
rect 2337 966 2343 1542
rect 2377 966 2383 1542
rect 2337 954 2383 966
rect 2455 1542 2501 1554
rect 2455 966 2461 1542
rect 2495 966 2501 1542
rect 2455 954 2501 966
rect 2573 1542 2619 1554
rect 2573 966 2579 1542
rect 2613 966 2619 1542
rect 2573 954 2619 966
rect 2691 1542 2737 1554
rect 2691 966 2697 1542
rect 2731 966 2737 1542
rect 2691 954 2737 966
rect 2809 1542 2855 1554
rect 2809 966 2815 1542
rect 2849 966 2855 1542
rect 2809 954 2855 966
rect 2927 1542 2973 1554
rect 2927 966 2933 1542
rect 2967 966 2973 1542
rect 2927 954 2973 966
rect -2920 907 -2862 913
rect -2920 873 -2908 907
rect -2874 873 -2862 907
rect -2920 867 -2862 873
rect -2802 907 -2744 913
rect -2802 873 -2790 907
rect -2756 873 -2744 907
rect -2802 867 -2744 873
rect -2684 907 -2626 913
rect -2684 873 -2672 907
rect -2638 873 -2626 907
rect -2684 867 -2626 873
rect -2566 907 -2508 913
rect -2566 873 -2554 907
rect -2520 873 -2508 907
rect -2566 867 -2508 873
rect -2448 907 -2390 913
rect -2448 873 -2436 907
rect -2402 873 -2390 907
rect -2448 867 -2390 873
rect -2330 907 -2272 913
rect -2330 873 -2318 907
rect -2284 873 -2272 907
rect -2330 867 -2272 873
rect -2212 907 -2154 913
rect -2212 873 -2200 907
rect -2166 873 -2154 907
rect -2212 867 -2154 873
rect -2094 907 -2036 913
rect -2094 873 -2082 907
rect -2048 873 -2036 907
rect -2094 867 -2036 873
rect -1976 907 -1918 913
rect -1976 873 -1964 907
rect -1930 873 -1918 907
rect -1976 867 -1918 873
rect -1858 907 -1800 913
rect -1858 873 -1846 907
rect -1812 873 -1800 907
rect -1858 867 -1800 873
rect -1740 907 -1682 913
rect -1740 873 -1728 907
rect -1694 873 -1682 907
rect -1740 867 -1682 873
rect -1622 907 -1564 913
rect -1622 873 -1610 907
rect -1576 873 -1564 907
rect -1622 867 -1564 873
rect -1504 907 -1446 913
rect -1504 873 -1492 907
rect -1458 873 -1446 907
rect -1504 867 -1446 873
rect -1386 907 -1328 913
rect -1386 873 -1374 907
rect -1340 873 -1328 907
rect -1386 867 -1328 873
rect -1268 907 -1210 913
rect -1268 873 -1256 907
rect -1222 873 -1210 907
rect -1268 867 -1210 873
rect -1150 907 -1092 913
rect -1150 873 -1138 907
rect -1104 873 -1092 907
rect -1150 867 -1092 873
rect -1032 907 -974 913
rect -1032 873 -1020 907
rect -986 873 -974 907
rect -1032 867 -974 873
rect -914 907 -856 913
rect -914 873 -902 907
rect -868 873 -856 907
rect -914 867 -856 873
rect -796 907 -738 913
rect -796 873 -784 907
rect -750 873 -738 907
rect -796 867 -738 873
rect -678 907 -620 913
rect -678 873 -666 907
rect -632 873 -620 907
rect -678 867 -620 873
rect -560 907 -502 913
rect -560 873 -548 907
rect -514 873 -502 907
rect -560 867 -502 873
rect -442 907 -384 913
rect -442 873 -430 907
rect -396 873 -384 907
rect -442 867 -384 873
rect -324 907 -266 913
rect -324 873 -312 907
rect -278 873 -266 907
rect -324 867 -266 873
rect -206 907 -148 913
rect -206 873 -194 907
rect -160 873 -148 907
rect -206 867 -148 873
rect -88 907 -30 913
rect -88 873 -76 907
rect -42 873 -30 907
rect -88 867 -30 873
rect 30 907 88 913
rect 30 873 42 907
rect 76 873 88 907
rect 30 867 88 873
rect 148 907 206 913
rect 148 873 160 907
rect 194 873 206 907
rect 148 867 206 873
rect 266 907 324 913
rect 266 873 278 907
rect 312 873 324 907
rect 266 867 324 873
rect 384 907 442 913
rect 384 873 396 907
rect 430 873 442 907
rect 384 867 442 873
rect 502 907 560 913
rect 502 873 514 907
rect 548 873 560 907
rect 502 867 560 873
rect 620 907 678 913
rect 620 873 632 907
rect 666 873 678 907
rect 620 867 678 873
rect 738 907 796 913
rect 738 873 750 907
rect 784 873 796 907
rect 738 867 796 873
rect 856 907 914 913
rect 856 873 868 907
rect 902 873 914 907
rect 856 867 914 873
rect 974 907 1032 913
rect 974 873 986 907
rect 1020 873 1032 907
rect 974 867 1032 873
rect 1092 907 1150 913
rect 1092 873 1104 907
rect 1138 873 1150 907
rect 1092 867 1150 873
rect 1210 907 1268 913
rect 1210 873 1222 907
rect 1256 873 1268 907
rect 1210 867 1268 873
rect 1328 907 1386 913
rect 1328 873 1340 907
rect 1374 873 1386 907
rect 1328 867 1386 873
rect 1446 907 1504 913
rect 1446 873 1458 907
rect 1492 873 1504 907
rect 1446 867 1504 873
rect 1564 907 1622 913
rect 1564 873 1576 907
rect 1610 873 1622 907
rect 1564 867 1622 873
rect 1682 907 1740 913
rect 1682 873 1694 907
rect 1728 873 1740 907
rect 1682 867 1740 873
rect 1800 907 1858 913
rect 1800 873 1812 907
rect 1846 873 1858 907
rect 1800 867 1858 873
rect 1918 907 1976 913
rect 1918 873 1930 907
rect 1964 873 1976 907
rect 1918 867 1976 873
rect 2036 907 2094 913
rect 2036 873 2048 907
rect 2082 873 2094 907
rect 2036 867 2094 873
rect 2154 907 2212 913
rect 2154 873 2166 907
rect 2200 873 2212 907
rect 2154 867 2212 873
rect 2272 907 2330 913
rect 2272 873 2284 907
rect 2318 873 2330 907
rect 2272 867 2330 873
rect 2390 907 2448 913
rect 2390 873 2402 907
rect 2436 873 2448 907
rect 2390 867 2448 873
rect 2508 907 2566 913
rect 2508 873 2520 907
rect 2554 873 2566 907
rect 2508 867 2566 873
rect 2626 907 2684 913
rect 2626 873 2638 907
rect 2672 873 2684 907
rect 2626 867 2684 873
rect 2744 907 2802 913
rect 2744 873 2756 907
rect 2790 873 2802 907
rect 2744 867 2802 873
rect 2862 907 2920 913
rect 2862 873 2874 907
rect 2908 873 2920 907
rect 2862 867 2920 873
rect -2920 799 -2862 805
rect -2920 765 -2908 799
rect -2874 765 -2862 799
rect -2920 759 -2862 765
rect -2802 799 -2744 805
rect -2802 765 -2790 799
rect -2756 765 -2744 799
rect -2802 759 -2744 765
rect -2684 799 -2626 805
rect -2684 765 -2672 799
rect -2638 765 -2626 799
rect -2684 759 -2626 765
rect -2566 799 -2508 805
rect -2566 765 -2554 799
rect -2520 765 -2508 799
rect -2566 759 -2508 765
rect -2448 799 -2390 805
rect -2448 765 -2436 799
rect -2402 765 -2390 799
rect -2448 759 -2390 765
rect -2330 799 -2272 805
rect -2330 765 -2318 799
rect -2284 765 -2272 799
rect -2330 759 -2272 765
rect -2212 799 -2154 805
rect -2212 765 -2200 799
rect -2166 765 -2154 799
rect -2212 759 -2154 765
rect -2094 799 -2036 805
rect -2094 765 -2082 799
rect -2048 765 -2036 799
rect -2094 759 -2036 765
rect -1976 799 -1918 805
rect -1976 765 -1964 799
rect -1930 765 -1918 799
rect -1976 759 -1918 765
rect -1858 799 -1800 805
rect -1858 765 -1846 799
rect -1812 765 -1800 799
rect -1858 759 -1800 765
rect -1740 799 -1682 805
rect -1740 765 -1728 799
rect -1694 765 -1682 799
rect -1740 759 -1682 765
rect -1622 799 -1564 805
rect -1622 765 -1610 799
rect -1576 765 -1564 799
rect -1622 759 -1564 765
rect -1504 799 -1446 805
rect -1504 765 -1492 799
rect -1458 765 -1446 799
rect -1504 759 -1446 765
rect -1386 799 -1328 805
rect -1386 765 -1374 799
rect -1340 765 -1328 799
rect -1386 759 -1328 765
rect -1268 799 -1210 805
rect -1268 765 -1256 799
rect -1222 765 -1210 799
rect -1268 759 -1210 765
rect -1150 799 -1092 805
rect -1150 765 -1138 799
rect -1104 765 -1092 799
rect -1150 759 -1092 765
rect -1032 799 -974 805
rect -1032 765 -1020 799
rect -986 765 -974 799
rect -1032 759 -974 765
rect -914 799 -856 805
rect -914 765 -902 799
rect -868 765 -856 799
rect -914 759 -856 765
rect -796 799 -738 805
rect -796 765 -784 799
rect -750 765 -738 799
rect -796 759 -738 765
rect -678 799 -620 805
rect -678 765 -666 799
rect -632 765 -620 799
rect -678 759 -620 765
rect -560 799 -502 805
rect -560 765 -548 799
rect -514 765 -502 799
rect -560 759 -502 765
rect -442 799 -384 805
rect -442 765 -430 799
rect -396 765 -384 799
rect -442 759 -384 765
rect -324 799 -266 805
rect -324 765 -312 799
rect -278 765 -266 799
rect -324 759 -266 765
rect -206 799 -148 805
rect -206 765 -194 799
rect -160 765 -148 799
rect -206 759 -148 765
rect -88 799 -30 805
rect -88 765 -76 799
rect -42 765 -30 799
rect -88 759 -30 765
rect 30 799 88 805
rect 30 765 42 799
rect 76 765 88 799
rect 30 759 88 765
rect 148 799 206 805
rect 148 765 160 799
rect 194 765 206 799
rect 148 759 206 765
rect 266 799 324 805
rect 266 765 278 799
rect 312 765 324 799
rect 266 759 324 765
rect 384 799 442 805
rect 384 765 396 799
rect 430 765 442 799
rect 384 759 442 765
rect 502 799 560 805
rect 502 765 514 799
rect 548 765 560 799
rect 502 759 560 765
rect 620 799 678 805
rect 620 765 632 799
rect 666 765 678 799
rect 620 759 678 765
rect 738 799 796 805
rect 738 765 750 799
rect 784 765 796 799
rect 738 759 796 765
rect 856 799 914 805
rect 856 765 868 799
rect 902 765 914 799
rect 856 759 914 765
rect 974 799 1032 805
rect 974 765 986 799
rect 1020 765 1032 799
rect 974 759 1032 765
rect 1092 799 1150 805
rect 1092 765 1104 799
rect 1138 765 1150 799
rect 1092 759 1150 765
rect 1210 799 1268 805
rect 1210 765 1222 799
rect 1256 765 1268 799
rect 1210 759 1268 765
rect 1328 799 1386 805
rect 1328 765 1340 799
rect 1374 765 1386 799
rect 1328 759 1386 765
rect 1446 799 1504 805
rect 1446 765 1458 799
rect 1492 765 1504 799
rect 1446 759 1504 765
rect 1564 799 1622 805
rect 1564 765 1576 799
rect 1610 765 1622 799
rect 1564 759 1622 765
rect 1682 799 1740 805
rect 1682 765 1694 799
rect 1728 765 1740 799
rect 1682 759 1740 765
rect 1800 799 1858 805
rect 1800 765 1812 799
rect 1846 765 1858 799
rect 1800 759 1858 765
rect 1918 799 1976 805
rect 1918 765 1930 799
rect 1964 765 1976 799
rect 1918 759 1976 765
rect 2036 799 2094 805
rect 2036 765 2048 799
rect 2082 765 2094 799
rect 2036 759 2094 765
rect 2154 799 2212 805
rect 2154 765 2166 799
rect 2200 765 2212 799
rect 2154 759 2212 765
rect 2272 799 2330 805
rect 2272 765 2284 799
rect 2318 765 2330 799
rect 2272 759 2330 765
rect 2390 799 2448 805
rect 2390 765 2402 799
rect 2436 765 2448 799
rect 2390 759 2448 765
rect 2508 799 2566 805
rect 2508 765 2520 799
rect 2554 765 2566 799
rect 2508 759 2566 765
rect 2626 799 2684 805
rect 2626 765 2638 799
rect 2672 765 2684 799
rect 2626 759 2684 765
rect 2744 799 2802 805
rect 2744 765 2756 799
rect 2790 765 2802 799
rect 2744 759 2802 765
rect 2862 799 2920 805
rect 2862 765 2874 799
rect 2908 765 2920 799
rect 2862 759 2920 765
rect -2973 706 -2927 718
rect -2973 130 -2967 706
rect -2933 130 -2927 706
rect -2973 118 -2927 130
rect -2855 706 -2809 718
rect -2855 130 -2849 706
rect -2815 130 -2809 706
rect -2855 118 -2809 130
rect -2737 706 -2691 718
rect -2737 130 -2731 706
rect -2697 130 -2691 706
rect -2737 118 -2691 130
rect -2619 706 -2573 718
rect -2619 130 -2613 706
rect -2579 130 -2573 706
rect -2619 118 -2573 130
rect -2501 706 -2455 718
rect -2501 130 -2495 706
rect -2461 130 -2455 706
rect -2501 118 -2455 130
rect -2383 706 -2337 718
rect -2383 130 -2377 706
rect -2343 130 -2337 706
rect -2383 118 -2337 130
rect -2265 706 -2219 718
rect -2265 130 -2259 706
rect -2225 130 -2219 706
rect -2265 118 -2219 130
rect -2147 706 -2101 718
rect -2147 130 -2141 706
rect -2107 130 -2101 706
rect -2147 118 -2101 130
rect -2029 706 -1983 718
rect -2029 130 -2023 706
rect -1989 130 -1983 706
rect -2029 118 -1983 130
rect -1911 706 -1865 718
rect -1911 130 -1905 706
rect -1871 130 -1865 706
rect -1911 118 -1865 130
rect -1793 706 -1747 718
rect -1793 130 -1787 706
rect -1753 130 -1747 706
rect -1793 118 -1747 130
rect -1675 706 -1629 718
rect -1675 130 -1669 706
rect -1635 130 -1629 706
rect -1675 118 -1629 130
rect -1557 706 -1511 718
rect -1557 130 -1551 706
rect -1517 130 -1511 706
rect -1557 118 -1511 130
rect -1439 706 -1393 718
rect -1439 130 -1433 706
rect -1399 130 -1393 706
rect -1439 118 -1393 130
rect -1321 706 -1275 718
rect -1321 130 -1315 706
rect -1281 130 -1275 706
rect -1321 118 -1275 130
rect -1203 706 -1157 718
rect -1203 130 -1197 706
rect -1163 130 -1157 706
rect -1203 118 -1157 130
rect -1085 706 -1039 718
rect -1085 130 -1079 706
rect -1045 130 -1039 706
rect -1085 118 -1039 130
rect -967 706 -921 718
rect -967 130 -961 706
rect -927 130 -921 706
rect -967 118 -921 130
rect -849 706 -803 718
rect -849 130 -843 706
rect -809 130 -803 706
rect -849 118 -803 130
rect -731 706 -685 718
rect -731 130 -725 706
rect -691 130 -685 706
rect -731 118 -685 130
rect -613 706 -567 718
rect -613 130 -607 706
rect -573 130 -567 706
rect -613 118 -567 130
rect -495 706 -449 718
rect -495 130 -489 706
rect -455 130 -449 706
rect -495 118 -449 130
rect -377 706 -331 718
rect -377 130 -371 706
rect -337 130 -331 706
rect -377 118 -331 130
rect -259 706 -213 718
rect -259 130 -253 706
rect -219 130 -213 706
rect -259 118 -213 130
rect -141 706 -95 718
rect -141 130 -135 706
rect -101 130 -95 706
rect -141 118 -95 130
rect -23 706 23 718
rect -23 130 -17 706
rect 17 130 23 706
rect -23 118 23 130
rect 95 706 141 718
rect 95 130 101 706
rect 135 130 141 706
rect 95 118 141 130
rect 213 706 259 718
rect 213 130 219 706
rect 253 130 259 706
rect 213 118 259 130
rect 331 706 377 718
rect 331 130 337 706
rect 371 130 377 706
rect 331 118 377 130
rect 449 706 495 718
rect 449 130 455 706
rect 489 130 495 706
rect 449 118 495 130
rect 567 706 613 718
rect 567 130 573 706
rect 607 130 613 706
rect 567 118 613 130
rect 685 706 731 718
rect 685 130 691 706
rect 725 130 731 706
rect 685 118 731 130
rect 803 706 849 718
rect 803 130 809 706
rect 843 130 849 706
rect 803 118 849 130
rect 921 706 967 718
rect 921 130 927 706
rect 961 130 967 706
rect 921 118 967 130
rect 1039 706 1085 718
rect 1039 130 1045 706
rect 1079 130 1085 706
rect 1039 118 1085 130
rect 1157 706 1203 718
rect 1157 130 1163 706
rect 1197 130 1203 706
rect 1157 118 1203 130
rect 1275 706 1321 718
rect 1275 130 1281 706
rect 1315 130 1321 706
rect 1275 118 1321 130
rect 1393 706 1439 718
rect 1393 130 1399 706
rect 1433 130 1439 706
rect 1393 118 1439 130
rect 1511 706 1557 718
rect 1511 130 1517 706
rect 1551 130 1557 706
rect 1511 118 1557 130
rect 1629 706 1675 718
rect 1629 130 1635 706
rect 1669 130 1675 706
rect 1629 118 1675 130
rect 1747 706 1793 718
rect 1747 130 1753 706
rect 1787 130 1793 706
rect 1747 118 1793 130
rect 1865 706 1911 718
rect 1865 130 1871 706
rect 1905 130 1911 706
rect 1865 118 1911 130
rect 1983 706 2029 718
rect 1983 130 1989 706
rect 2023 130 2029 706
rect 1983 118 2029 130
rect 2101 706 2147 718
rect 2101 130 2107 706
rect 2141 130 2147 706
rect 2101 118 2147 130
rect 2219 706 2265 718
rect 2219 130 2225 706
rect 2259 130 2265 706
rect 2219 118 2265 130
rect 2337 706 2383 718
rect 2337 130 2343 706
rect 2377 130 2383 706
rect 2337 118 2383 130
rect 2455 706 2501 718
rect 2455 130 2461 706
rect 2495 130 2501 706
rect 2455 118 2501 130
rect 2573 706 2619 718
rect 2573 130 2579 706
rect 2613 130 2619 706
rect 2573 118 2619 130
rect 2691 706 2737 718
rect 2691 130 2697 706
rect 2731 130 2737 706
rect 2691 118 2737 130
rect 2809 706 2855 718
rect 2809 130 2815 706
rect 2849 130 2855 706
rect 2809 118 2855 130
rect 2927 706 2973 718
rect 2927 130 2933 706
rect 2967 130 2973 706
rect 2927 118 2973 130
rect -2920 71 -2862 77
rect -2920 37 -2908 71
rect -2874 37 -2862 71
rect -2920 31 -2862 37
rect -2802 71 -2744 77
rect -2802 37 -2790 71
rect -2756 37 -2744 71
rect -2802 31 -2744 37
rect -2684 71 -2626 77
rect -2684 37 -2672 71
rect -2638 37 -2626 71
rect -2684 31 -2626 37
rect -2566 71 -2508 77
rect -2566 37 -2554 71
rect -2520 37 -2508 71
rect -2566 31 -2508 37
rect -2448 71 -2390 77
rect -2448 37 -2436 71
rect -2402 37 -2390 71
rect -2448 31 -2390 37
rect -2330 71 -2272 77
rect -2330 37 -2318 71
rect -2284 37 -2272 71
rect -2330 31 -2272 37
rect -2212 71 -2154 77
rect -2212 37 -2200 71
rect -2166 37 -2154 71
rect -2212 31 -2154 37
rect -2094 71 -2036 77
rect -2094 37 -2082 71
rect -2048 37 -2036 71
rect -2094 31 -2036 37
rect -1976 71 -1918 77
rect -1976 37 -1964 71
rect -1930 37 -1918 71
rect -1976 31 -1918 37
rect -1858 71 -1800 77
rect -1858 37 -1846 71
rect -1812 37 -1800 71
rect -1858 31 -1800 37
rect -1740 71 -1682 77
rect -1740 37 -1728 71
rect -1694 37 -1682 71
rect -1740 31 -1682 37
rect -1622 71 -1564 77
rect -1622 37 -1610 71
rect -1576 37 -1564 71
rect -1622 31 -1564 37
rect -1504 71 -1446 77
rect -1504 37 -1492 71
rect -1458 37 -1446 71
rect -1504 31 -1446 37
rect -1386 71 -1328 77
rect -1386 37 -1374 71
rect -1340 37 -1328 71
rect -1386 31 -1328 37
rect -1268 71 -1210 77
rect -1268 37 -1256 71
rect -1222 37 -1210 71
rect -1268 31 -1210 37
rect -1150 71 -1092 77
rect -1150 37 -1138 71
rect -1104 37 -1092 71
rect -1150 31 -1092 37
rect -1032 71 -974 77
rect -1032 37 -1020 71
rect -986 37 -974 71
rect -1032 31 -974 37
rect -914 71 -856 77
rect -914 37 -902 71
rect -868 37 -856 71
rect -914 31 -856 37
rect -796 71 -738 77
rect -796 37 -784 71
rect -750 37 -738 71
rect -796 31 -738 37
rect -678 71 -620 77
rect -678 37 -666 71
rect -632 37 -620 71
rect -678 31 -620 37
rect -560 71 -502 77
rect -560 37 -548 71
rect -514 37 -502 71
rect -560 31 -502 37
rect -442 71 -384 77
rect -442 37 -430 71
rect -396 37 -384 71
rect -442 31 -384 37
rect -324 71 -266 77
rect -324 37 -312 71
rect -278 37 -266 71
rect -324 31 -266 37
rect -206 71 -148 77
rect -206 37 -194 71
rect -160 37 -148 71
rect -206 31 -148 37
rect -88 71 -30 77
rect -88 37 -76 71
rect -42 37 -30 71
rect -88 31 -30 37
rect 30 71 88 77
rect 30 37 42 71
rect 76 37 88 71
rect 30 31 88 37
rect 148 71 206 77
rect 148 37 160 71
rect 194 37 206 71
rect 148 31 206 37
rect 266 71 324 77
rect 266 37 278 71
rect 312 37 324 71
rect 266 31 324 37
rect 384 71 442 77
rect 384 37 396 71
rect 430 37 442 71
rect 384 31 442 37
rect 502 71 560 77
rect 502 37 514 71
rect 548 37 560 71
rect 502 31 560 37
rect 620 71 678 77
rect 620 37 632 71
rect 666 37 678 71
rect 620 31 678 37
rect 738 71 796 77
rect 738 37 750 71
rect 784 37 796 71
rect 738 31 796 37
rect 856 71 914 77
rect 856 37 868 71
rect 902 37 914 71
rect 856 31 914 37
rect 974 71 1032 77
rect 974 37 986 71
rect 1020 37 1032 71
rect 974 31 1032 37
rect 1092 71 1150 77
rect 1092 37 1104 71
rect 1138 37 1150 71
rect 1092 31 1150 37
rect 1210 71 1268 77
rect 1210 37 1222 71
rect 1256 37 1268 71
rect 1210 31 1268 37
rect 1328 71 1386 77
rect 1328 37 1340 71
rect 1374 37 1386 71
rect 1328 31 1386 37
rect 1446 71 1504 77
rect 1446 37 1458 71
rect 1492 37 1504 71
rect 1446 31 1504 37
rect 1564 71 1622 77
rect 1564 37 1576 71
rect 1610 37 1622 71
rect 1564 31 1622 37
rect 1682 71 1740 77
rect 1682 37 1694 71
rect 1728 37 1740 71
rect 1682 31 1740 37
rect 1800 71 1858 77
rect 1800 37 1812 71
rect 1846 37 1858 71
rect 1800 31 1858 37
rect 1918 71 1976 77
rect 1918 37 1930 71
rect 1964 37 1976 71
rect 1918 31 1976 37
rect 2036 71 2094 77
rect 2036 37 2048 71
rect 2082 37 2094 71
rect 2036 31 2094 37
rect 2154 71 2212 77
rect 2154 37 2166 71
rect 2200 37 2212 71
rect 2154 31 2212 37
rect 2272 71 2330 77
rect 2272 37 2284 71
rect 2318 37 2330 71
rect 2272 31 2330 37
rect 2390 71 2448 77
rect 2390 37 2402 71
rect 2436 37 2448 71
rect 2390 31 2448 37
rect 2508 71 2566 77
rect 2508 37 2520 71
rect 2554 37 2566 71
rect 2508 31 2566 37
rect 2626 71 2684 77
rect 2626 37 2638 71
rect 2672 37 2684 71
rect 2626 31 2684 37
rect 2744 71 2802 77
rect 2744 37 2756 71
rect 2790 37 2802 71
rect 2744 31 2802 37
rect 2862 71 2920 77
rect 2862 37 2874 71
rect 2908 37 2920 71
rect 2862 31 2920 37
rect -2920 -37 -2862 -31
rect -2920 -71 -2908 -37
rect -2874 -71 -2862 -37
rect -2920 -77 -2862 -71
rect -2802 -37 -2744 -31
rect -2802 -71 -2790 -37
rect -2756 -71 -2744 -37
rect -2802 -77 -2744 -71
rect -2684 -37 -2626 -31
rect -2684 -71 -2672 -37
rect -2638 -71 -2626 -37
rect -2684 -77 -2626 -71
rect -2566 -37 -2508 -31
rect -2566 -71 -2554 -37
rect -2520 -71 -2508 -37
rect -2566 -77 -2508 -71
rect -2448 -37 -2390 -31
rect -2448 -71 -2436 -37
rect -2402 -71 -2390 -37
rect -2448 -77 -2390 -71
rect -2330 -37 -2272 -31
rect -2330 -71 -2318 -37
rect -2284 -71 -2272 -37
rect -2330 -77 -2272 -71
rect -2212 -37 -2154 -31
rect -2212 -71 -2200 -37
rect -2166 -71 -2154 -37
rect -2212 -77 -2154 -71
rect -2094 -37 -2036 -31
rect -2094 -71 -2082 -37
rect -2048 -71 -2036 -37
rect -2094 -77 -2036 -71
rect -1976 -37 -1918 -31
rect -1976 -71 -1964 -37
rect -1930 -71 -1918 -37
rect -1976 -77 -1918 -71
rect -1858 -37 -1800 -31
rect -1858 -71 -1846 -37
rect -1812 -71 -1800 -37
rect -1858 -77 -1800 -71
rect -1740 -37 -1682 -31
rect -1740 -71 -1728 -37
rect -1694 -71 -1682 -37
rect -1740 -77 -1682 -71
rect -1622 -37 -1564 -31
rect -1622 -71 -1610 -37
rect -1576 -71 -1564 -37
rect -1622 -77 -1564 -71
rect -1504 -37 -1446 -31
rect -1504 -71 -1492 -37
rect -1458 -71 -1446 -37
rect -1504 -77 -1446 -71
rect -1386 -37 -1328 -31
rect -1386 -71 -1374 -37
rect -1340 -71 -1328 -37
rect -1386 -77 -1328 -71
rect -1268 -37 -1210 -31
rect -1268 -71 -1256 -37
rect -1222 -71 -1210 -37
rect -1268 -77 -1210 -71
rect -1150 -37 -1092 -31
rect -1150 -71 -1138 -37
rect -1104 -71 -1092 -37
rect -1150 -77 -1092 -71
rect -1032 -37 -974 -31
rect -1032 -71 -1020 -37
rect -986 -71 -974 -37
rect -1032 -77 -974 -71
rect -914 -37 -856 -31
rect -914 -71 -902 -37
rect -868 -71 -856 -37
rect -914 -77 -856 -71
rect -796 -37 -738 -31
rect -796 -71 -784 -37
rect -750 -71 -738 -37
rect -796 -77 -738 -71
rect -678 -37 -620 -31
rect -678 -71 -666 -37
rect -632 -71 -620 -37
rect -678 -77 -620 -71
rect -560 -37 -502 -31
rect -560 -71 -548 -37
rect -514 -71 -502 -37
rect -560 -77 -502 -71
rect -442 -37 -384 -31
rect -442 -71 -430 -37
rect -396 -71 -384 -37
rect -442 -77 -384 -71
rect -324 -37 -266 -31
rect -324 -71 -312 -37
rect -278 -71 -266 -37
rect -324 -77 -266 -71
rect -206 -37 -148 -31
rect -206 -71 -194 -37
rect -160 -71 -148 -37
rect -206 -77 -148 -71
rect -88 -37 -30 -31
rect -88 -71 -76 -37
rect -42 -71 -30 -37
rect -88 -77 -30 -71
rect 30 -37 88 -31
rect 30 -71 42 -37
rect 76 -71 88 -37
rect 30 -77 88 -71
rect 148 -37 206 -31
rect 148 -71 160 -37
rect 194 -71 206 -37
rect 148 -77 206 -71
rect 266 -37 324 -31
rect 266 -71 278 -37
rect 312 -71 324 -37
rect 266 -77 324 -71
rect 384 -37 442 -31
rect 384 -71 396 -37
rect 430 -71 442 -37
rect 384 -77 442 -71
rect 502 -37 560 -31
rect 502 -71 514 -37
rect 548 -71 560 -37
rect 502 -77 560 -71
rect 620 -37 678 -31
rect 620 -71 632 -37
rect 666 -71 678 -37
rect 620 -77 678 -71
rect 738 -37 796 -31
rect 738 -71 750 -37
rect 784 -71 796 -37
rect 738 -77 796 -71
rect 856 -37 914 -31
rect 856 -71 868 -37
rect 902 -71 914 -37
rect 856 -77 914 -71
rect 974 -37 1032 -31
rect 974 -71 986 -37
rect 1020 -71 1032 -37
rect 974 -77 1032 -71
rect 1092 -37 1150 -31
rect 1092 -71 1104 -37
rect 1138 -71 1150 -37
rect 1092 -77 1150 -71
rect 1210 -37 1268 -31
rect 1210 -71 1222 -37
rect 1256 -71 1268 -37
rect 1210 -77 1268 -71
rect 1328 -37 1386 -31
rect 1328 -71 1340 -37
rect 1374 -71 1386 -37
rect 1328 -77 1386 -71
rect 1446 -37 1504 -31
rect 1446 -71 1458 -37
rect 1492 -71 1504 -37
rect 1446 -77 1504 -71
rect 1564 -37 1622 -31
rect 1564 -71 1576 -37
rect 1610 -71 1622 -37
rect 1564 -77 1622 -71
rect 1682 -37 1740 -31
rect 1682 -71 1694 -37
rect 1728 -71 1740 -37
rect 1682 -77 1740 -71
rect 1800 -37 1858 -31
rect 1800 -71 1812 -37
rect 1846 -71 1858 -37
rect 1800 -77 1858 -71
rect 1918 -37 1976 -31
rect 1918 -71 1930 -37
rect 1964 -71 1976 -37
rect 1918 -77 1976 -71
rect 2036 -37 2094 -31
rect 2036 -71 2048 -37
rect 2082 -71 2094 -37
rect 2036 -77 2094 -71
rect 2154 -37 2212 -31
rect 2154 -71 2166 -37
rect 2200 -71 2212 -37
rect 2154 -77 2212 -71
rect 2272 -37 2330 -31
rect 2272 -71 2284 -37
rect 2318 -71 2330 -37
rect 2272 -77 2330 -71
rect 2390 -37 2448 -31
rect 2390 -71 2402 -37
rect 2436 -71 2448 -37
rect 2390 -77 2448 -71
rect 2508 -37 2566 -31
rect 2508 -71 2520 -37
rect 2554 -71 2566 -37
rect 2508 -77 2566 -71
rect 2626 -37 2684 -31
rect 2626 -71 2638 -37
rect 2672 -71 2684 -37
rect 2626 -77 2684 -71
rect 2744 -37 2802 -31
rect 2744 -71 2756 -37
rect 2790 -71 2802 -37
rect 2744 -77 2802 -71
rect 2862 -37 2920 -31
rect 2862 -71 2874 -37
rect 2908 -71 2920 -37
rect 2862 -77 2920 -71
rect -2973 -130 -2927 -118
rect -2973 -706 -2967 -130
rect -2933 -706 -2927 -130
rect -2973 -718 -2927 -706
rect -2855 -130 -2809 -118
rect -2855 -706 -2849 -130
rect -2815 -706 -2809 -130
rect -2855 -718 -2809 -706
rect -2737 -130 -2691 -118
rect -2737 -706 -2731 -130
rect -2697 -706 -2691 -130
rect -2737 -718 -2691 -706
rect -2619 -130 -2573 -118
rect -2619 -706 -2613 -130
rect -2579 -706 -2573 -130
rect -2619 -718 -2573 -706
rect -2501 -130 -2455 -118
rect -2501 -706 -2495 -130
rect -2461 -706 -2455 -130
rect -2501 -718 -2455 -706
rect -2383 -130 -2337 -118
rect -2383 -706 -2377 -130
rect -2343 -706 -2337 -130
rect -2383 -718 -2337 -706
rect -2265 -130 -2219 -118
rect -2265 -706 -2259 -130
rect -2225 -706 -2219 -130
rect -2265 -718 -2219 -706
rect -2147 -130 -2101 -118
rect -2147 -706 -2141 -130
rect -2107 -706 -2101 -130
rect -2147 -718 -2101 -706
rect -2029 -130 -1983 -118
rect -2029 -706 -2023 -130
rect -1989 -706 -1983 -130
rect -2029 -718 -1983 -706
rect -1911 -130 -1865 -118
rect -1911 -706 -1905 -130
rect -1871 -706 -1865 -130
rect -1911 -718 -1865 -706
rect -1793 -130 -1747 -118
rect -1793 -706 -1787 -130
rect -1753 -706 -1747 -130
rect -1793 -718 -1747 -706
rect -1675 -130 -1629 -118
rect -1675 -706 -1669 -130
rect -1635 -706 -1629 -130
rect -1675 -718 -1629 -706
rect -1557 -130 -1511 -118
rect -1557 -706 -1551 -130
rect -1517 -706 -1511 -130
rect -1557 -718 -1511 -706
rect -1439 -130 -1393 -118
rect -1439 -706 -1433 -130
rect -1399 -706 -1393 -130
rect -1439 -718 -1393 -706
rect -1321 -130 -1275 -118
rect -1321 -706 -1315 -130
rect -1281 -706 -1275 -130
rect -1321 -718 -1275 -706
rect -1203 -130 -1157 -118
rect -1203 -706 -1197 -130
rect -1163 -706 -1157 -130
rect -1203 -718 -1157 -706
rect -1085 -130 -1039 -118
rect -1085 -706 -1079 -130
rect -1045 -706 -1039 -130
rect -1085 -718 -1039 -706
rect -967 -130 -921 -118
rect -967 -706 -961 -130
rect -927 -706 -921 -130
rect -967 -718 -921 -706
rect -849 -130 -803 -118
rect -849 -706 -843 -130
rect -809 -706 -803 -130
rect -849 -718 -803 -706
rect -731 -130 -685 -118
rect -731 -706 -725 -130
rect -691 -706 -685 -130
rect -731 -718 -685 -706
rect -613 -130 -567 -118
rect -613 -706 -607 -130
rect -573 -706 -567 -130
rect -613 -718 -567 -706
rect -495 -130 -449 -118
rect -495 -706 -489 -130
rect -455 -706 -449 -130
rect -495 -718 -449 -706
rect -377 -130 -331 -118
rect -377 -706 -371 -130
rect -337 -706 -331 -130
rect -377 -718 -331 -706
rect -259 -130 -213 -118
rect -259 -706 -253 -130
rect -219 -706 -213 -130
rect -259 -718 -213 -706
rect -141 -130 -95 -118
rect -141 -706 -135 -130
rect -101 -706 -95 -130
rect -141 -718 -95 -706
rect -23 -130 23 -118
rect -23 -706 -17 -130
rect 17 -706 23 -130
rect -23 -718 23 -706
rect 95 -130 141 -118
rect 95 -706 101 -130
rect 135 -706 141 -130
rect 95 -718 141 -706
rect 213 -130 259 -118
rect 213 -706 219 -130
rect 253 -706 259 -130
rect 213 -718 259 -706
rect 331 -130 377 -118
rect 331 -706 337 -130
rect 371 -706 377 -130
rect 331 -718 377 -706
rect 449 -130 495 -118
rect 449 -706 455 -130
rect 489 -706 495 -130
rect 449 -718 495 -706
rect 567 -130 613 -118
rect 567 -706 573 -130
rect 607 -706 613 -130
rect 567 -718 613 -706
rect 685 -130 731 -118
rect 685 -706 691 -130
rect 725 -706 731 -130
rect 685 -718 731 -706
rect 803 -130 849 -118
rect 803 -706 809 -130
rect 843 -706 849 -130
rect 803 -718 849 -706
rect 921 -130 967 -118
rect 921 -706 927 -130
rect 961 -706 967 -130
rect 921 -718 967 -706
rect 1039 -130 1085 -118
rect 1039 -706 1045 -130
rect 1079 -706 1085 -130
rect 1039 -718 1085 -706
rect 1157 -130 1203 -118
rect 1157 -706 1163 -130
rect 1197 -706 1203 -130
rect 1157 -718 1203 -706
rect 1275 -130 1321 -118
rect 1275 -706 1281 -130
rect 1315 -706 1321 -130
rect 1275 -718 1321 -706
rect 1393 -130 1439 -118
rect 1393 -706 1399 -130
rect 1433 -706 1439 -130
rect 1393 -718 1439 -706
rect 1511 -130 1557 -118
rect 1511 -706 1517 -130
rect 1551 -706 1557 -130
rect 1511 -718 1557 -706
rect 1629 -130 1675 -118
rect 1629 -706 1635 -130
rect 1669 -706 1675 -130
rect 1629 -718 1675 -706
rect 1747 -130 1793 -118
rect 1747 -706 1753 -130
rect 1787 -706 1793 -130
rect 1747 -718 1793 -706
rect 1865 -130 1911 -118
rect 1865 -706 1871 -130
rect 1905 -706 1911 -130
rect 1865 -718 1911 -706
rect 1983 -130 2029 -118
rect 1983 -706 1989 -130
rect 2023 -706 2029 -130
rect 1983 -718 2029 -706
rect 2101 -130 2147 -118
rect 2101 -706 2107 -130
rect 2141 -706 2147 -130
rect 2101 -718 2147 -706
rect 2219 -130 2265 -118
rect 2219 -706 2225 -130
rect 2259 -706 2265 -130
rect 2219 -718 2265 -706
rect 2337 -130 2383 -118
rect 2337 -706 2343 -130
rect 2377 -706 2383 -130
rect 2337 -718 2383 -706
rect 2455 -130 2501 -118
rect 2455 -706 2461 -130
rect 2495 -706 2501 -130
rect 2455 -718 2501 -706
rect 2573 -130 2619 -118
rect 2573 -706 2579 -130
rect 2613 -706 2619 -130
rect 2573 -718 2619 -706
rect 2691 -130 2737 -118
rect 2691 -706 2697 -130
rect 2731 -706 2737 -130
rect 2691 -718 2737 -706
rect 2809 -130 2855 -118
rect 2809 -706 2815 -130
rect 2849 -706 2855 -130
rect 2809 -718 2855 -706
rect 2927 -130 2973 -118
rect 2927 -706 2933 -130
rect 2967 -706 2973 -130
rect 2927 -718 2973 -706
rect -2920 -765 -2862 -759
rect -2920 -799 -2908 -765
rect -2874 -799 -2862 -765
rect -2920 -805 -2862 -799
rect -2802 -765 -2744 -759
rect -2802 -799 -2790 -765
rect -2756 -799 -2744 -765
rect -2802 -805 -2744 -799
rect -2684 -765 -2626 -759
rect -2684 -799 -2672 -765
rect -2638 -799 -2626 -765
rect -2684 -805 -2626 -799
rect -2566 -765 -2508 -759
rect -2566 -799 -2554 -765
rect -2520 -799 -2508 -765
rect -2566 -805 -2508 -799
rect -2448 -765 -2390 -759
rect -2448 -799 -2436 -765
rect -2402 -799 -2390 -765
rect -2448 -805 -2390 -799
rect -2330 -765 -2272 -759
rect -2330 -799 -2318 -765
rect -2284 -799 -2272 -765
rect -2330 -805 -2272 -799
rect -2212 -765 -2154 -759
rect -2212 -799 -2200 -765
rect -2166 -799 -2154 -765
rect -2212 -805 -2154 -799
rect -2094 -765 -2036 -759
rect -2094 -799 -2082 -765
rect -2048 -799 -2036 -765
rect -2094 -805 -2036 -799
rect -1976 -765 -1918 -759
rect -1976 -799 -1964 -765
rect -1930 -799 -1918 -765
rect -1976 -805 -1918 -799
rect -1858 -765 -1800 -759
rect -1858 -799 -1846 -765
rect -1812 -799 -1800 -765
rect -1858 -805 -1800 -799
rect -1740 -765 -1682 -759
rect -1740 -799 -1728 -765
rect -1694 -799 -1682 -765
rect -1740 -805 -1682 -799
rect -1622 -765 -1564 -759
rect -1622 -799 -1610 -765
rect -1576 -799 -1564 -765
rect -1622 -805 -1564 -799
rect -1504 -765 -1446 -759
rect -1504 -799 -1492 -765
rect -1458 -799 -1446 -765
rect -1504 -805 -1446 -799
rect -1386 -765 -1328 -759
rect -1386 -799 -1374 -765
rect -1340 -799 -1328 -765
rect -1386 -805 -1328 -799
rect -1268 -765 -1210 -759
rect -1268 -799 -1256 -765
rect -1222 -799 -1210 -765
rect -1268 -805 -1210 -799
rect -1150 -765 -1092 -759
rect -1150 -799 -1138 -765
rect -1104 -799 -1092 -765
rect -1150 -805 -1092 -799
rect -1032 -765 -974 -759
rect -1032 -799 -1020 -765
rect -986 -799 -974 -765
rect -1032 -805 -974 -799
rect -914 -765 -856 -759
rect -914 -799 -902 -765
rect -868 -799 -856 -765
rect -914 -805 -856 -799
rect -796 -765 -738 -759
rect -796 -799 -784 -765
rect -750 -799 -738 -765
rect -796 -805 -738 -799
rect -678 -765 -620 -759
rect -678 -799 -666 -765
rect -632 -799 -620 -765
rect -678 -805 -620 -799
rect -560 -765 -502 -759
rect -560 -799 -548 -765
rect -514 -799 -502 -765
rect -560 -805 -502 -799
rect -442 -765 -384 -759
rect -442 -799 -430 -765
rect -396 -799 -384 -765
rect -442 -805 -384 -799
rect -324 -765 -266 -759
rect -324 -799 -312 -765
rect -278 -799 -266 -765
rect -324 -805 -266 -799
rect -206 -765 -148 -759
rect -206 -799 -194 -765
rect -160 -799 -148 -765
rect -206 -805 -148 -799
rect -88 -765 -30 -759
rect -88 -799 -76 -765
rect -42 -799 -30 -765
rect -88 -805 -30 -799
rect 30 -765 88 -759
rect 30 -799 42 -765
rect 76 -799 88 -765
rect 30 -805 88 -799
rect 148 -765 206 -759
rect 148 -799 160 -765
rect 194 -799 206 -765
rect 148 -805 206 -799
rect 266 -765 324 -759
rect 266 -799 278 -765
rect 312 -799 324 -765
rect 266 -805 324 -799
rect 384 -765 442 -759
rect 384 -799 396 -765
rect 430 -799 442 -765
rect 384 -805 442 -799
rect 502 -765 560 -759
rect 502 -799 514 -765
rect 548 -799 560 -765
rect 502 -805 560 -799
rect 620 -765 678 -759
rect 620 -799 632 -765
rect 666 -799 678 -765
rect 620 -805 678 -799
rect 738 -765 796 -759
rect 738 -799 750 -765
rect 784 -799 796 -765
rect 738 -805 796 -799
rect 856 -765 914 -759
rect 856 -799 868 -765
rect 902 -799 914 -765
rect 856 -805 914 -799
rect 974 -765 1032 -759
rect 974 -799 986 -765
rect 1020 -799 1032 -765
rect 974 -805 1032 -799
rect 1092 -765 1150 -759
rect 1092 -799 1104 -765
rect 1138 -799 1150 -765
rect 1092 -805 1150 -799
rect 1210 -765 1268 -759
rect 1210 -799 1222 -765
rect 1256 -799 1268 -765
rect 1210 -805 1268 -799
rect 1328 -765 1386 -759
rect 1328 -799 1340 -765
rect 1374 -799 1386 -765
rect 1328 -805 1386 -799
rect 1446 -765 1504 -759
rect 1446 -799 1458 -765
rect 1492 -799 1504 -765
rect 1446 -805 1504 -799
rect 1564 -765 1622 -759
rect 1564 -799 1576 -765
rect 1610 -799 1622 -765
rect 1564 -805 1622 -799
rect 1682 -765 1740 -759
rect 1682 -799 1694 -765
rect 1728 -799 1740 -765
rect 1682 -805 1740 -799
rect 1800 -765 1858 -759
rect 1800 -799 1812 -765
rect 1846 -799 1858 -765
rect 1800 -805 1858 -799
rect 1918 -765 1976 -759
rect 1918 -799 1930 -765
rect 1964 -799 1976 -765
rect 1918 -805 1976 -799
rect 2036 -765 2094 -759
rect 2036 -799 2048 -765
rect 2082 -799 2094 -765
rect 2036 -805 2094 -799
rect 2154 -765 2212 -759
rect 2154 -799 2166 -765
rect 2200 -799 2212 -765
rect 2154 -805 2212 -799
rect 2272 -765 2330 -759
rect 2272 -799 2284 -765
rect 2318 -799 2330 -765
rect 2272 -805 2330 -799
rect 2390 -765 2448 -759
rect 2390 -799 2402 -765
rect 2436 -799 2448 -765
rect 2390 -805 2448 -799
rect 2508 -765 2566 -759
rect 2508 -799 2520 -765
rect 2554 -799 2566 -765
rect 2508 -805 2566 -799
rect 2626 -765 2684 -759
rect 2626 -799 2638 -765
rect 2672 -799 2684 -765
rect 2626 -805 2684 -799
rect 2744 -765 2802 -759
rect 2744 -799 2756 -765
rect 2790 -799 2802 -765
rect 2744 -805 2802 -799
rect 2862 -765 2920 -759
rect 2862 -799 2874 -765
rect 2908 -799 2920 -765
rect 2862 -805 2920 -799
rect -2920 -873 -2862 -867
rect -2920 -907 -2908 -873
rect -2874 -907 -2862 -873
rect -2920 -913 -2862 -907
rect -2802 -873 -2744 -867
rect -2802 -907 -2790 -873
rect -2756 -907 -2744 -873
rect -2802 -913 -2744 -907
rect -2684 -873 -2626 -867
rect -2684 -907 -2672 -873
rect -2638 -907 -2626 -873
rect -2684 -913 -2626 -907
rect -2566 -873 -2508 -867
rect -2566 -907 -2554 -873
rect -2520 -907 -2508 -873
rect -2566 -913 -2508 -907
rect -2448 -873 -2390 -867
rect -2448 -907 -2436 -873
rect -2402 -907 -2390 -873
rect -2448 -913 -2390 -907
rect -2330 -873 -2272 -867
rect -2330 -907 -2318 -873
rect -2284 -907 -2272 -873
rect -2330 -913 -2272 -907
rect -2212 -873 -2154 -867
rect -2212 -907 -2200 -873
rect -2166 -907 -2154 -873
rect -2212 -913 -2154 -907
rect -2094 -873 -2036 -867
rect -2094 -907 -2082 -873
rect -2048 -907 -2036 -873
rect -2094 -913 -2036 -907
rect -1976 -873 -1918 -867
rect -1976 -907 -1964 -873
rect -1930 -907 -1918 -873
rect -1976 -913 -1918 -907
rect -1858 -873 -1800 -867
rect -1858 -907 -1846 -873
rect -1812 -907 -1800 -873
rect -1858 -913 -1800 -907
rect -1740 -873 -1682 -867
rect -1740 -907 -1728 -873
rect -1694 -907 -1682 -873
rect -1740 -913 -1682 -907
rect -1622 -873 -1564 -867
rect -1622 -907 -1610 -873
rect -1576 -907 -1564 -873
rect -1622 -913 -1564 -907
rect -1504 -873 -1446 -867
rect -1504 -907 -1492 -873
rect -1458 -907 -1446 -873
rect -1504 -913 -1446 -907
rect -1386 -873 -1328 -867
rect -1386 -907 -1374 -873
rect -1340 -907 -1328 -873
rect -1386 -913 -1328 -907
rect -1268 -873 -1210 -867
rect -1268 -907 -1256 -873
rect -1222 -907 -1210 -873
rect -1268 -913 -1210 -907
rect -1150 -873 -1092 -867
rect -1150 -907 -1138 -873
rect -1104 -907 -1092 -873
rect -1150 -913 -1092 -907
rect -1032 -873 -974 -867
rect -1032 -907 -1020 -873
rect -986 -907 -974 -873
rect -1032 -913 -974 -907
rect -914 -873 -856 -867
rect -914 -907 -902 -873
rect -868 -907 -856 -873
rect -914 -913 -856 -907
rect -796 -873 -738 -867
rect -796 -907 -784 -873
rect -750 -907 -738 -873
rect -796 -913 -738 -907
rect -678 -873 -620 -867
rect -678 -907 -666 -873
rect -632 -907 -620 -873
rect -678 -913 -620 -907
rect -560 -873 -502 -867
rect -560 -907 -548 -873
rect -514 -907 -502 -873
rect -560 -913 -502 -907
rect -442 -873 -384 -867
rect -442 -907 -430 -873
rect -396 -907 -384 -873
rect -442 -913 -384 -907
rect -324 -873 -266 -867
rect -324 -907 -312 -873
rect -278 -907 -266 -873
rect -324 -913 -266 -907
rect -206 -873 -148 -867
rect -206 -907 -194 -873
rect -160 -907 -148 -873
rect -206 -913 -148 -907
rect -88 -873 -30 -867
rect -88 -907 -76 -873
rect -42 -907 -30 -873
rect -88 -913 -30 -907
rect 30 -873 88 -867
rect 30 -907 42 -873
rect 76 -907 88 -873
rect 30 -913 88 -907
rect 148 -873 206 -867
rect 148 -907 160 -873
rect 194 -907 206 -873
rect 148 -913 206 -907
rect 266 -873 324 -867
rect 266 -907 278 -873
rect 312 -907 324 -873
rect 266 -913 324 -907
rect 384 -873 442 -867
rect 384 -907 396 -873
rect 430 -907 442 -873
rect 384 -913 442 -907
rect 502 -873 560 -867
rect 502 -907 514 -873
rect 548 -907 560 -873
rect 502 -913 560 -907
rect 620 -873 678 -867
rect 620 -907 632 -873
rect 666 -907 678 -873
rect 620 -913 678 -907
rect 738 -873 796 -867
rect 738 -907 750 -873
rect 784 -907 796 -873
rect 738 -913 796 -907
rect 856 -873 914 -867
rect 856 -907 868 -873
rect 902 -907 914 -873
rect 856 -913 914 -907
rect 974 -873 1032 -867
rect 974 -907 986 -873
rect 1020 -907 1032 -873
rect 974 -913 1032 -907
rect 1092 -873 1150 -867
rect 1092 -907 1104 -873
rect 1138 -907 1150 -873
rect 1092 -913 1150 -907
rect 1210 -873 1268 -867
rect 1210 -907 1222 -873
rect 1256 -907 1268 -873
rect 1210 -913 1268 -907
rect 1328 -873 1386 -867
rect 1328 -907 1340 -873
rect 1374 -907 1386 -873
rect 1328 -913 1386 -907
rect 1446 -873 1504 -867
rect 1446 -907 1458 -873
rect 1492 -907 1504 -873
rect 1446 -913 1504 -907
rect 1564 -873 1622 -867
rect 1564 -907 1576 -873
rect 1610 -907 1622 -873
rect 1564 -913 1622 -907
rect 1682 -873 1740 -867
rect 1682 -907 1694 -873
rect 1728 -907 1740 -873
rect 1682 -913 1740 -907
rect 1800 -873 1858 -867
rect 1800 -907 1812 -873
rect 1846 -907 1858 -873
rect 1800 -913 1858 -907
rect 1918 -873 1976 -867
rect 1918 -907 1930 -873
rect 1964 -907 1976 -873
rect 1918 -913 1976 -907
rect 2036 -873 2094 -867
rect 2036 -907 2048 -873
rect 2082 -907 2094 -873
rect 2036 -913 2094 -907
rect 2154 -873 2212 -867
rect 2154 -907 2166 -873
rect 2200 -907 2212 -873
rect 2154 -913 2212 -907
rect 2272 -873 2330 -867
rect 2272 -907 2284 -873
rect 2318 -907 2330 -873
rect 2272 -913 2330 -907
rect 2390 -873 2448 -867
rect 2390 -907 2402 -873
rect 2436 -907 2448 -873
rect 2390 -913 2448 -907
rect 2508 -873 2566 -867
rect 2508 -907 2520 -873
rect 2554 -907 2566 -873
rect 2508 -913 2566 -907
rect 2626 -873 2684 -867
rect 2626 -907 2638 -873
rect 2672 -907 2684 -873
rect 2626 -913 2684 -907
rect 2744 -873 2802 -867
rect 2744 -907 2756 -873
rect 2790 -907 2802 -873
rect 2744 -913 2802 -907
rect 2862 -873 2920 -867
rect 2862 -907 2874 -873
rect 2908 -907 2920 -873
rect 2862 -913 2920 -907
rect -2973 -966 -2927 -954
rect -2973 -1542 -2967 -966
rect -2933 -1542 -2927 -966
rect -2973 -1554 -2927 -1542
rect -2855 -966 -2809 -954
rect -2855 -1542 -2849 -966
rect -2815 -1542 -2809 -966
rect -2855 -1554 -2809 -1542
rect -2737 -966 -2691 -954
rect -2737 -1542 -2731 -966
rect -2697 -1542 -2691 -966
rect -2737 -1554 -2691 -1542
rect -2619 -966 -2573 -954
rect -2619 -1542 -2613 -966
rect -2579 -1542 -2573 -966
rect -2619 -1554 -2573 -1542
rect -2501 -966 -2455 -954
rect -2501 -1542 -2495 -966
rect -2461 -1542 -2455 -966
rect -2501 -1554 -2455 -1542
rect -2383 -966 -2337 -954
rect -2383 -1542 -2377 -966
rect -2343 -1542 -2337 -966
rect -2383 -1554 -2337 -1542
rect -2265 -966 -2219 -954
rect -2265 -1542 -2259 -966
rect -2225 -1542 -2219 -966
rect -2265 -1554 -2219 -1542
rect -2147 -966 -2101 -954
rect -2147 -1542 -2141 -966
rect -2107 -1542 -2101 -966
rect -2147 -1554 -2101 -1542
rect -2029 -966 -1983 -954
rect -2029 -1542 -2023 -966
rect -1989 -1542 -1983 -966
rect -2029 -1554 -1983 -1542
rect -1911 -966 -1865 -954
rect -1911 -1542 -1905 -966
rect -1871 -1542 -1865 -966
rect -1911 -1554 -1865 -1542
rect -1793 -966 -1747 -954
rect -1793 -1542 -1787 -966
rect -1753 -1542 -1747 -966
rect -1793 -1554 -1747 -1542
rect -1675 -966 -1629 -954
rect -1675 -1542 -1669 -966
rect -1635 -1542 -1629 -966
rect -1675 -1554 -1629 -1542
rect -1557 -966 -1511 -954
rect -1557 -1542 -1551 -966
rect -1517 -1542 -1511 -966
rect -1557 -1554 -1511 -1542
rect -1439 -966 -1393 -954
rect -1439 -1542 -1433 -966
rect -1399 -1542 -1393 -966
rect -1439 -1554 -1393 -1542
rect -1321 -966 -1275 -954
rect -1321 -1542 -1315 -966
rect -1281 -1542 -1275 -966
rect -1321 -1554 -1275 -1542
rect -1203 -966 -1157 -954
rect -1203 -1542 -1197 -966
rect -1163 -1542 -1157 -966
rect -1203 -1554 -1157 -1542
rect -1085 -966 -1039 -954
rect -1085 -1542 -1079 -966
rect -1045 -1542 -1039 -966
rect -1085 -1554 -1039 -1542
rect -967 -966 -921 -954
rect -967 -1542 -961 -966
rect -927 -1542 -921 -966
rect -967 -1554 -921 -1542
rect -849 -966 -803 -954
rect -849 -1542 -843 -966
rect -809 -1542 -803 -966
rect -849 -1554 -803 -1542
rect -731 -966 -685 -954
rect -731 -1542 -725 -966
rect -691 -1542 -685 -966
rect -731 -1554 -685 -1542
rect -613 -966 -567 -954
rect -613 -1542 -607 -966
rect -573 -1542 -567 -966
rect -613 -1554 -567 -1542
rect -495 -966 -449 -954
rect -495 -1542 -489 -966
rect -455 -1542 -449 -966
rect -495 -1554 -449 -1542
rect -377 -966 -331 -954
rect -377 -1542 -371 -966
rect -337 -1542 -331 -966
rect -377 -1554 -331 -1542
rect -259 -966 -213 -954
rect -259 -1542 -253 -966
rect -219 -1542 -213 -966
rect -259 -1554 -213 -1542
rect -141 -966 -95 -954
rect -141 -1542 -135 -966
rect -101 -1542 -95 -966
rect -141 -1554 -95 -1542
rect -23 -966 23 -954
rect -23 -1542 -17 -966
rect 17 -1542 23 -966
rect -23 -1554 23 -1542
rect 95 -966 141 -954
rect 95 -1542 101 -966
rect 135 -1542 141 -966
rect 95 -1554 141 -1542
rect 213 -966 259 -954
rect 213 -1542 219 -966
rect 253 -1542 259 -966
rect 213 -1554 259 -1542
rect 331 -966 377 -954
rect 331 -1542 337 -966
rect 371 -1542 377 -966
rect 331 -1554 377 -1542
rect 449 -966 495 -954
rect 449 -1542 455 -966
rect 489 -1542 495 -966
rect 449 -1554 495 -1542
rect 567 -966 613 -954
rect 567 -1542 573 -966
rect 607 -1542 613 -966
rect 567 -1554 613 -1542
rect 685 -966 731 -954
rect 685 -1542 691 -966
rect 725 -1542 731 -966
rect 685 -1554 731 -1542
rect 803 -966 849 -954
rect 803 -1542 809 -966
rect 843 -1542 849 -966
rect 803 -1554 849 -1542
rect 921 -966 967 -954
rect 921 -1542 927 -966
rect 961 -1542 967 -966
rect 921 -1554 967 -1542
rect 1039 -966 1085 -954
rect 1039 -1542 1045 -966
rect 1079 -1542 1085 -966
rect 1039 -1554 1085 -1542
rect 1157 -966 1203 -954
rect 1157 -1542 1163 -966
rect 1197 -1542 1203 -966
rect 1157 -1554 1203 -1542
rect 1275 -966 1321 -954
rect 1275 -1542 1281 -966
rect 1315 -1542 1321 -966
rect 1275 -1554 1321 -1542
rect 1393 -966 1439 -954
rect 1393 -1542 1399 -966
rect 1433 -1542 1439 -966
rect 1393 -1554 1439 -1542
rect 1511 -966 1557 -954
rect 1511 -1542 1517 -966
rect 1551 -1542 1557 -966
rect 1511 -1554 1557 -1542
rect 1629 -966 1675 -954
rect 1629 -1542 1635 -966
rect 1669 -1542 1675 -966
rect 1629 -1554 1675 -1542
rect 1747 -966 1793 -954
rect 1747 -1542 1753 -966
rect 1787 -1542 1793 -966
rect 1747 -1554 1793 -1542
rect 1865 -966 1911 -954
rect 1865 -1542 1871 -966
rect 1905 -1542 1911 -966
rect 1865 -1554 1911 -1542
rect 1983 -966 2029 -954
rect 1983 -1542 1989 -966
rect 2023 -1542 2029 -966
rect 1983 -1554 2029 -1542
rect 2101 -966 2147 -954
rect 2101 -1542 2107 -966
rect 2141 -1542 2147 -966
rect 2101 -1554 2147 -1542
rect 2219 -966 2265 -954
rect 2219 -1542 2225 -966
rect 2259 -1542 2265 -966
rect 2219 -1554 2265 -1542
rect 2337 -966 2383 -954
rect 2337 -1542 2343 -966
rect 2377 -1542 2383 -966
rect 2337 -1554 2383 -1542
rect 2455 -966 2501 -954
rect 2455 -1542 2461 -966
rect 2495 -1542 2501 -966
rect 2455 -1554 2501 -1542
rect 2573 -966 2619 -954
rect 2573 -1542 2579 -966
rect 2613 -1542 2619 -966
rect 2573 -1554 2619 -1542
rect 2691 -966 2737 -954
rect 2691 -1542 2697 -966
rect 2731 -1542 2737 -966
rect 2691 -1554 2737 -1542
rect 2809 -966 2855 -954
rect 2809 -1542 2815 -966
rect 2849 -1542 2855 -966
rect 2809 -1554 2855 -1542
rect 2927 -966 2973 -954
rect 2927 -1542 2933 -966
rect 2967 -1542 2973 -966
rect 2927 -1554 2973 -1542
rect -2920 -1601 -2862 -1595
rect -2920 -1635 -2908 -1601
rect -2874 -1635 -2862 -1601
rect -2920 -1641 -2862 -1635
rect -2802 -1601 -2744 -1595
rect -2802 -1635 -2790 -1601
rect -2756 -1635 -2744 -1601
rect -2802 -1641 -2744 -1635
rect -2684 -1601 -2626 -1595
rect -2684 -1635 -2672 -1601
rect -2638 -1635 -2626 -1601
rect -2684 -1641 -2626 -1635
rect -2566 -1601 -2508 -1595
rect -2566 -1635 -2554 -1601
rect -2520 -1635 -2508 -1601
rect -2566 -1641 -2508 -1635
rect -2448 -1601 -2390 -1595
rect -2448 -1635 -2436 -1601
rect -2402 -1635 -2390 -1601
rect -2448 -1641 -2390 -1635
rect -2330 -1601 -2272 -1595
rect -2330 -1635 -2318 -1601
rect -2284 -1635 -2272 -1601
rect -2330 -1641 -2272 -1635
rect -2212 -1601 -2154 -1595
rect -2212 -1635 -2200 -1601
rect -2166 -1635 -2154 -1601
rect -2212 -1641 -2154 -1635
rect -2094 -1601 -2036 -1595
rect -2094 -1635 -2082 -1601
rect -2048 -1635 -2036 -1601
rect -2094 -1641 -2036 -1635
rect -1976 -1601 -1918 -1595
rect -1976 -1635 -1964 -1601
rect -1930 -1635 -1918 -1601
rect -1976 -1641 -1918 -1635
rect -1858 -1601 -1800 -1595
rect -1858 -1635 -1846 -1601
rect -1812 -1635 -1800 -1601
rect -1858 -1641 -1800 -1635
rect -1740 -1601 -1682 -1595
rect -1740 -1635 -1728 -1601
rect -1694 -1635 -1682 -1601
rect -1740 -1641 -1682 -1635
rect -1622 -1601 -1564 -1595
rect -1622 -1635 -1610 -1601
rect -1576 -1635 -1564 -1601
rect -1622 -1641 -1564 -1635
rect -1504 -1601 -1446 -1595
rect -1504 -1635 -1492 -1601
rect -1458 -1635 -1446 -1601
rect -1504 -1641 -1446 -1635
rect -1386 -1601 -1328 -1595
rect -1386 -1635 -1374 -1601
rect -1340 -1635 -1328 -1601
rect -1386 -1641 -1328 -1635
rect -1268 -1601 -1210 -1595
rect -1268 -1635 -1256 -1601
rect -1222 -1635 -1210 -1601
rect -1268 -1641 -1210 -1635
rect -1150 -1601 -1092 -1595
rect -1150 -1635 -1138 -1601
rect -1104 -1635 -1092 -1601
rect -1150 -1641 -1092 -1635
rect -1032 -1601 -974 -1595
rect -1032 -1635 -1020 -1601
rect -986 -1635 -974 -1601
rect -1032 -1641 -974 -1635
rect -914 -1601 -856 -1595
rect -914 -1635 -902 -1601
rect -868 -1635 -856 -1601
rect -914 -1641 -856 -1635
rect -796 -1601 -738 -1595
rect -796 -1635 -784 -1601
rect -750 -1635 -738 -1601
rect -796 -1641 -738 -1635
rect -678 -1601 -620 -1595
rect -678 -1635 -666 -1601
rect -632 -1635 -620 -1601
rect -678 -1641 -620 -1635
rect -560 -1601 -502 -1595
rect -560 -1635 -548 -1601
rect -514 -1635 -502 -1601
rect -560 -1641 -502 -1635
rect -442 -1601 -384 -1595
rect -442 -1635 -430 -1601
rect -396 -1635 -384 -1601
rect -442 -1641 -384 -1635
rect -324 -1601 -266 -1595
rect -324 -1635 -312 -1601
rect -278 -1635 -266 -1601
rect -324 -1641 -266 -1635
rect -206 -1601 -148 -1595
rect -206 -1635 -194 -1601
rect -160 -1635 -148 -1601
rect -206 -1641 -148 -1635
rect -88 -1601 -30 -1595
rect -88 -1635 -76 -1601
rect -42 -1635 -30 -1601
rect -88 -1641 -30 -1635
rect 30 -1601 88 -1595
rect 30 -1635 42 -1601
rect 76 -1635 88 -1601
rect 30 -1641 88 -1635
rect 148 -1601 206 -1595
rect 148 -1635 160 -1601
rect 194 -1635 206 -1601
rect 148 -1641 206 -1635
rect 266 -1601 324 -1595
rect 266 -1635 278 -1601
rect 312 -1635 324 -1601
rect 266 -1641 324 -1635
rect 384 -1601 442 -1595
rect 384 -1635 396 -1601
rect 430 -1635 442 -1601
rect 384 -1641 442 -1635
rect 502 -1601 560 -1595
rect 502 -1635 514 -1601
rect 548 -1635 560 -1601
rect 502 -1641 560 -1635
rect 620 -1601 678 -1595
rect 620 -1635 632 -1601
rect 666 -1635 678 -1601
rect 620 -1641 678 -1635
rect 738 -1601 796 -1595
rect 738 -1635 750 -1601
rect 784 -1635 796 -1601
rect 738 -1641 796 -1635
rect 856 -1601 914 -1595
rect 856 -1635 868 -1601
rect 902 -1635 914 -1601
rect 856 -1641 914 -1635
rect 974 -1601 1032 -1595
rect 974 -1635 986 -1601
rect 1020 -1635 1032 -1601
rect 974 -1641 1032 -1635
rect 1092 -1601 1150 -1595
rect 1092 -1635 1104 -1601
rect 1138 -1635 1150 -1601
rect 1092 -1641 1150 -1635
rect 1210 -1601 1268 -1595
rect 1210 -1635 1222 -1601
rect 1256 -1635 1268 -1601
rect 1210 -1641 1268 -1635
rect 1328 -1601 1386 -1595
rect 1328 -1635 1340 -1601
rect 1374 -1635 1386 -1601
rect 1328 -1641 1386 -1635
rect 1446 -1601 1504 -1595
rect 1446 -1635 1458 -1601
rect 1492 -1635 1504 -1601
rect 1446 -1641 1504 -1635
rect 1564 -1601 1622 -1595
rect 1564 -1635 1576 -1601
rect 1610 -1635 1622 -1601
rect 1564 -1641 1622 -1635
rect 1682 -1601 1740 -1595
rect 1682 -1635 1694 -1601
rect 1728 -1635 1740 -1601
rect 1682 -1641 1740 -1635
rect 1800 -1601 1858 -1595
rect 1800 -1635 1812 -1601
rect 1846 -1635 1858 -1601
rect 1800 -1641 1858 -1635
rect 1918 -1601 1976 -1595
rect 1918 -1635 1930 -1601
rect 1964 -1635 1976 -1601
rect 1918 -1641 1976 -1635
rect 2036 -1601 2094 -1595
rect 2036 -1635 2048 -1601
rect 2082 -1635 2094 -1601
rect 2036 -1641 2094 -1635
rect 2154 -1601 2212 -1595
rect 2154 -1635 2166 -1601
rect 2200 -1635 2212 -1601
rect 2154 -1641 2212 -1635
rect 2272 -1601 2330 -1595
rect 2272 -1635 2284 -1601
rect 2318 -1635 2330 -1601
rect 2272 -1641 2330 -1635
rect 2390 -1601 2448 -1595
rect 2390 -1635 2402 -1601
rect 2436 -1635 2448 -1601
rect 2390 -1641 2448 -1635
rect 2508 -1601 2566 -1595
rect 2508 -1635 2520 -1601
rect 2554 -1635 2566 -1601
rect 2508 -1641 2566 -1635
rect 2626 -1601 2684 -1595
rect 2626 -1635 2638 -1601
rect 2672 -1635 2684 -1601
rect 2626 -1641 2684 -1635
rect 2744 -1601 2802 -1595
rect 2744 -1635 2756 -1601
rect 2790 -1635 2802 -1601
rect 2744 -1641 2802 -1635
rect 2862 -1601 2920 -1595
rect 2862 -1635 2874 -1601
rect 2908 -1635 2920 -1601
rect 2862 -1641 2920 -1635
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -3064 -1720 3064 1720
string parameters w 3 l 0.3 m 4 nf 50 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
