magic
tech sky130B
magscale 1 2
timestamp 1606423877
<< error_p >>
rect -2920 1217 -2862 1223
rect -2802 1217 -2744 1223
rect -2684 1217 -2626 1223
rect -2566 1217 -2508 1223
rect -2448 1217 -2390 1223
rect -2330 1217 -2272 1223
rect -2212 1217 -2154 1223
rect -2094 1217 -2036 1223
rect -1976 1217 -1918 1223
rect -1858 1217 -1800 1223
rect -1740 1217 -1682 1223
rect -1622 1217 -1564 1223
rect -1504 1217 -1446 1223
rect -1386 1217 -1328 1223
rect -1268 1217 -1210 1223
rect -1150 1217 -1092 1223
rect -1032 1217 -974 1223
rect -914 1217 -856 1223
rect -796 1217 -738 1223
rect -678 1217 -620 1223
rect -560 1217 -502 1223
rect -442 1217 -384 1223
rect -324 1217 -266 1223
rect -206 1217 -148 1223
rect -88 1217 -30 1223
rect 30 1217 88 1223
rect 148 1217 206 1223
rect 266 1217 324 1223
rect 384 1217 442 1223
rect 502 1217 560 1223
rect 620 1217 678 1223
rect 738 1217 796 1223
rect 856 1217 914 1223
rect 974 1217 1032 1223
rect 1092 1217 1150 1223
rect 1210 1217 1268 1223
rect 1328 1217 1386 1223
rect 1446 1217 1504 1223
rect 1564 1217 1622 1223
rect 1682 1217 1740 1223
rect 1800 1217 1858 1223
rect 1918 1217 1976 1223
rect 2036 1217 2094 1223
rect 2154 1217 2212 1223
rect 2272 1217 2330 1223
rect 2390 1217 2448 1223
rect 2508 1217 2566 1223
rect 2626 1217 2684 1223
rect 2744 1217 2802 1223
rect 2862 1217 2920 1223
rect -2920 1183 -2908 1217
rect -2802 1183 -2790 1217
rect -2684 1183 -2672 1217
rect -2566 1183 -2554 1217
rect -2448 1183 -2436 1217
rect -2330 1183 -2318 1217
rect -2212 1183 -2200 1217
rect -2094 1183 -2082 1217
rect -1976 1183 -1964 1217
rect -1858 1183 -1846 1217
rect -1740 1183 -1728 1217
rect -1622 1183 -1610 1217
rect -1504 1183 -1492 1217
rect -1386 1183 -1374 1217
rect -1268 1183 -1256 1217
rect -1150 1183 -1138 1217
rect -1032 1183 -1020 1217
rect -914 1183 -902 1217
rect -796 1183 -784 1217
rect -678 1183 -666 1217
rect -560 1183 -548 1217
rect -442 1183 -430 1217
rect -324 1183 -312 1217
rect -206 1183 -194 1217
rect -88 1183 -76 1217
rect 30 1183 42 1217
rect 148 1183 160 1217
rect 266 1183 278 1217
rect 384 1183 396 1217
rect 502 1183 514 1217
rect 620 1183 632 1217
rect 738 1183 750 1217
rect 856 1183 868 1217
rect 974 1183 986 1217
rect 1092 1183 1104 1217
rect 1210 1183 1222 1217
rect 1328 1183 1340 1217
rect 1446 1183 1458 1217
rect 1564 1183 1576 1217
rect 1682 1183 1694 1217
rect 1800 1183 1812 1217
rect 1918 1183 1930 1217
rect 2036 1183 2048 1217
rect 2154 1183 2166 1217
rect 2272 1183 2284 1217
rect 2390 1183 2402 1217
rect 2508 1183 2520 1217
rect 2626 1183 2638 1217
rect 2744 1183 2756 1217
rect 2862 1183 2874 1217
rect -2920 1177 -2862 1183
rect -2802 1177 -2744 1183
rect -2684 1177 -2626 1183
rect -2566 1177 -2508 1183
rect -2448 1177 -2390 1183
rect -2330 1177 -2272 1183
rect -2212 1177 -2154 1183
rect -2094 1177 -2036 1183
rect -1976 1177 -1918 1183
rect -1858 1177 -1800 1183
rect -1740 1177 -1682 1183
rect -1622 1177 -1564 1183
rect -1504 1177 -1446 1183
rect -1386 1177 -1328 1183
rect -1268 1177 -1210 1183
rect -1150 1177 -1092 1183
rect -1032 1177 -974 1183
rect -914 1177 -856 1183
rect -796 1177 -738 1183
rect -678 1177 -620 1183
rect -560 1177 -502 1183
rect -442 1177 -384 1183
rect -324 1177 -266 1183
rect -206 1177 -148 1183
rect -88 1177 -30 1183
rect 30 1177 88 1183
rect 148 1177 206 1183
rect 266 1177 324 1183
rect 384 1177 442 1183
rect 502 1177 560 1183
rect 620 1177 678 1183
rect 738 1177 796 1183
rect 856 1177 914 1183
rect 974 1177 1032 1183
rect 1092 1177 1150 1183
rect 1210 1177 1268 1183
rect 1328 1177 1386 1183
rect 1446 1177 1504 1183
rect 1564 1177 1622 1183
rect 1682 1177 1740 1183
rect 1800 1177 1858 1183
rect 1918 1177 1976 1183
rect 2036 1177 2094 1183
rect 2154 1177 2212 1183
rect 2272 1177 2330 1183
rect 2390 1177 2448 1183
rect 2508 1177 2566 1183
rect 2626 1177 2684 1183
rect 2744 1177 2802 1183
rect 2862 1177 2920 1183
rect -2920 489 -2862 495
rect -2802 489 -2744 495
rect -2684 489 -2626 495
rect -2566 489 -2508 495
rect -2448 489 -2390 495
rect -2330 489 -2272 495
rect -2212 489 -2154 495
rect -2094 489 -2036 495
rect -1976 489 -1918 495
rect -1858 489 -1800 495
rect -1740 489 -1682 495
rect -1622 489 -1564 495
rect -1504 489 -1446 495
rect -1386 489 -1328 495
rect -1268 489 -1210 495
rect -1150 489 -1092 495
rect -1032 489 -974 495
rect -914 489 -856 495
rect -796 489 -738 495
rect -678 489 -620 495
rect -560 489 -502 495
rect -442 489 -384 495
rect -324 489 -266 495
rect -206 489 -148 495
rect -88 489 -30 495
rect 30 489 88 495
rect 148 489 206 495
rect 266 489 324 495
rect 384 489 442 495
rect 502 489 560 495
rect 620 489 678 495
rect 738 489 796 495
rect 856 489 914 495
rect 974 489 1032 495
rect 1092 489 1150 495
rect 1210 489 1268 495
rect 1328 489 1386 495
rect 1446 489 1504 495
rect 1564 489 1622 495
rect 1682 489 1740 495
rect 1800 489 1858 495
rect 1918 489 1976 495
rect 2036 489 2094 495
rect 2154 489 2212 495
rect 2272 489 2330 495
rect 2390 489 2448 495
rect 2508 489 2566 495
rect 2626 489 2684 495
rect 2744 489 2802 495
rect 2862 489 2920 495
rect -2920 455 -2908 489
rect -2802 455 -2790 489
rect -2684 455 -2672 489
rect -2566 455 -2554 489
rect -2448 455 -2436 489
rect -2330 455 -2318 489
rect -2212 455 -2200 489
rect -2094 455 -2082 489
rect -1976 455 -1964 489
rect -1858 455 -1846 489
rect -1740 455 -1728 489
rect -1622 455 -1610 489
rect -1504 455 -1492 489
rect -1386 455 -1374 489
rect -1268 455 -1256 489
rect -1150 455 -1138 489
rect -1032 455 -1020 489
rect -914 455 -902 489
rect -796 455 -784 489
rect -678 455 -666 489
rect -560 455 -548 489
rect -442 455 -430 489
rect -324 455 -312 489
rect -206 455 -194 489
rect -88 455 -76 489
rect 30 455 42 489
rect 148 455 160 489
rect 266 455 278 489
rect 384 455 396 489
rect 502 455 514 489
rect 620 455 632 489
rect 738 455 750 489
rect 856 455 868 489
rect 974 455 986 489
rect 1092 455 1104 489
rect 1210 455 1222 489
rect 1328 455 1340 489
rect 1446 455 1458 489
rect 1564 455 1576 489
rect 1682 455 1694 489
rect 1800 455 1812 489
rect 1918 455 1930 489
rect 2036 455 2048 489
rect 2154 455 2166 489
rect 2272 455 2284 489
rect 2390 455 2402 489
rect 2508 455 2520 489
rect 2626 455 2638 489
rect 2744 455 2756 489
rect 2862 455 2874 489
rect -2920 449 -2862 455
rect -2802 449 -2744 455
rect -2684 449 -2626 455
rect -2566 449 -2508 455
rect -2448 449 -2390 455
rect -2330 449 -2272 455
rect -2212 449 -2154 455
rect -2094 449 -2036 455
rect -1976 449 -1918 455
rect -1858 449 -1800 455
rect -1740 449 -1682 455
rect -1622 449 -1564 455
rect -1504 449 -1446 455
rect -1386 449 -1328 455
rect -1268 449 -1210 455
rect -1150 449 -1092 455
rect -1032 449 -974 455
rect -914 449 -856 455
rect -796 449 -738 455
rect -678 449 -620 455
rect -560 449 -502 455
rect -442 449 -384 455
rect -324 449 -266 455
rect -206 449 -148 455
rect -88 449 -30 455
rect 30 449 88 455
rect 148 449 206 455
rect 266 449 324 455
rect 384 449 442 455
rect 502 449 560 455
rect 620 449 678 455
rect 738 449 796 455
rect 856 449 914 455
rect 974 449 1032 455
rect 1092 449 1150 455
rect 1210 449 1268 455
rect 1328 449 1386 455
rect 1446 449 1504 455
rect 1564 449 1622 455
rect 1682 449 1740 455
rect 1800 449 1858 455
rect 1918 449 1976 455
rect 2036 449 2094 455
rect 2154 449 2212 455
rect 2272 449 2330 455
rect 2390 449 2448 455
rect 2508 449 2566 455
rect 2626 449 2684 455
rect 2744 449 2802 455
rect 2862 449 2920 455
rect -2920 381 -2862 387
rect -2802 381 -2744 387
rect -2684 381 -2626 387
rect -2566 381 -2508 387
rect -2448 381 -2390 387
rect -2330 381 -2272 387
rect -2212 381 -2154 387
rect -2094 381 -2036 387
rect -1976 381 -1918 387
rect -1858 381 -1800 387
rect -1740 381 -1682 387
rect -1622 381 -1564 387
rect -1504 381 -1446 387
rect -1386 381 -1328 387
rect -1268 381 -1210 387
rect -1150 381 -1092 387
rect -1032 381 -974 387
rect -914 381 -856 387
rect -796 381 -738 387
rect -678 381 -620 387
rect -560 381 -502 387
rect -442 381 -384 387
rect -324 381 -266 387
rect -206 381 -148 387
rect -88 381 -30 387
rect 30 381 88 387
rect 148 381 206 387
rect 266 381 324 387
rect 384 381 442 387
rect 502 381 560 387
rect 620 381 678 387
rect 738 381 796 387
rect 856 381 914 387
rect 974 381 1032 387
rect 1092 381 1150 387
rect 1210 381 1268 387
rect 1328 381 1386 387
rect 1446 381 1504 387
rect 1564 381 1622 387
rect 1682 381 1740 387
rect 1800 381 1858 387
rect 1918 381 1976 387
rect 2036 381 2094 387
rect 2154 381 2212 387
rect 2272 381 2330 387
rect 2390 381 2448 387
rect 2508 381 2566 387
rect 2626 381 2684 387
rect 2744 381 2802 387
rect 2862 381 2920 387
rect -2920 347 -2908 381
rect -2802 347 -2790 381
rect -2684 347 -2672 381
rect -2566 347 -2554 381
rect -2448 347 -2436 381
rect -2330 347 -2318 381
rect -2212 347 -2200 381
rect -2094 347 -2082 381
rect -1976 347 -1964 381
rect -1858 347 -1846 381
rect -1740 347 -1728 381
rect -1622 347 -1610 381
rect -1504 347 -1492 381
rect -1386 347 -1374 381
rect -1268 347 -1256 381
rect -1150 347 -1138 381
rect -1032 347 -1020 381
rect -914 347 -902 381
rect -796 347 -784 381
rect -678 347 -666 381
rect -560 347 -548 381
rect -442 347 -430 381
rect -324 347 -312 381
rect -206 347 -194 381
rect -88 347 -76 381
rect 30 347 42 381
rect 148 347 160 381
rect 266 347 278 381
rect 384 347 396 381
rect 502 347 514 381
rect 620 347 632 381
rect 738 347 750 381
rect 856 347 868 381
rect 974 347 986 381
rect 1092 347 1104 381
rect 1210 347 1222 381
rect 1328 347 1340 381
rect 1446 347 1458 381
rect 1564 347 1576 381
rect 1682 347 1694 381
rect 1800 347 1812 381
rect 1918 347 1930 381
rect 2036 347 2048 381
rect 2154 347 2166 381
rect 2272 347 2284 381
rect 2390 347 2402 381
rect 2508 347 2520 381
rect 2626 347 2638 381
rect 2744 347 2756 381
rect 2862 347 2874 381
rect -2920 341 -2862 347
rect -2802 341 -2744 347
rect -2684 341 -2626 347
rect -2566 341 -2508 347
rect -2448 341 -2390 347
rect -2330 341 -2272 347
rect -2212 341 -2154 347
rect -2094 341 -2036 347
rect -1976 341 -1918 347
rect -1858 341 -1800 347
rect -1740 341 -1682 347
rect -1622 341 -1564 347
rect -1504 341 -1446 347
rect -1386 341 -1328 347
rect -1268 341 -1210 347
rect -1150 341 -1092 347
rect -1032 341 -974 347
rect -914 341 -856 347
rect -796 341 -738 347
rect -678 341 -620 347
rect -560 341 -502 347
rect -442 341 -384 347
rect -324 341 -266 347
rect -206 341 -148 347
rect -88 341 -30 347
rect 30 341 88 347
rect 148 341 206 347
rect 266 341 324 347
rect 384 341 442 347
rect 502 341 560 347
rect 620 341 678 347
rect 738 341 796 347
rect 856 341 914 347
rect 974 341 1032 347
rect 1092 341 1150 347
rect 1210 341 1268 347
rect 1328 341 1386 347
rect 1446 341 1504 347
rect 1564 341 1622 347
rect 1682 341 1740 347
rect 1800 341 1858 347
rect 1918 341 1976 347
rect 2036 341 2094 347
rect 2154 341 2212 347
rect 2272 341 2330 347
rect 2390 341 2448 347
rect 2508 341 2566 347
rect 2626 341 2684 347
rect 2744 341 2802 347
rect 2862 341 2920 347
rect -2920 -347 -2862 -341
rect -2802 -347 -2744 -341
rect -2684 -347 -2626 -341
rect -2566 -347 -2508 -341
rect -2448 -347 -2390 -341
rect -2330 -347 -2272 -341
rect -2212 -347 -2154 -341
rect -2094 -347 -2036 -341
rect -1976 -347 -1918 -341
rect -1858 -347 -1800 -341
rect -1740 -347 -1682 -341
rect -1622 -347 -1564 -341
rect -1504 -347 -1446 -341
rect -1386 -347 -1328 -341
rect -1268 -347 -1210 -341
rect -1150 -347 -1092 -341
rect -1032 -347 -974 -341
rect -914 -347 -856 -341
rect -796 -347 -738 -341
rect -678 -347 -620 -341
rect -560 -347 -502 -341
rect -442 -347 -384 -341
rect -324 -347 -266 -341
rect -206 -347 -148 -341
rect -88 -347 -30 -341
rect 30 -347 88 -341
rect 148 -347 206 -341
rect 266 -347 324 -341
rect 384 -347 442 -341
rect 502 -347 560 -341
rect 620 -347 678 -341
rect 738 -347 796 -341
rect 856 -347 914 -341
rect 974 -347 1032 -341
rect 1092 -347 1150 -341
rect 1210 -347 1268 -341
rect 1328 -347 1386 -341
rect 1446 -347 1504 -341
rect 1564 -347 1622 -341
rect 1682 -347 1740 -341
rect 1800 -347 1858 -341
rect 1918 -347 1976 -341
rect 2036 -347 2094 -341
rect 2154 -347 2212 -341
rect 2272 -347 2330 -341
rect 2390 -347 2448 -341
rect 2508 -347 2566 -341
rect 2626 -347 2684 -341
rect 2744 -347 2802 -341
rect 2862 -347 2920 -341
rect -2920 -381 -2908 -347
rect -2802 -381 -2790 -347
rect -2684 -381 -2672 -347
rect -2566 -381 -2554 -347
rect -2448 -381 -2436 -347
rect -2330 -381 -2318 -347
rect -2212 -381 -2200 -347
rect -2094 -381 -2082 -347
rect -1976 -381 -1964 -347
rect -1858 -381 -1846 -347
rect -1740 -381 -1728 -347
rect -1622 -381 -1610 -347
rect -1504 -381 -1492 -347
rect -1386 -381 -1374 -347
rect -1268 -381 -1256 -347
rect -1150 -381 -1138 -347
rect -1032 -381 -1020 -347
rect -914 -381 -902 -347
rect -796 -381 -784 -347
rect -678 -381 -666 -347
rect -560 -381 -548 -347
rect -442 -381 -430 -347
rect -324 -381 -312 -347
rect -206 -381 -194 -347
rect -88 -381 -76 -347
rect 30 -381 42 -347
rect 148 -381 160 -347
rect 266 -381 278 -347
rect 384 -381 396 -347
rect 502 -381 514 -347
rect 620 -381 632 -347
rect 738 -381 750 -347
rect 856 -381 868 -347
rect 974 -381 986 -347
rect 1092 -381 1104 -347
rect 1210 -381 1222 -347
rect 1328 -381 1340 -347
rect 1446 -381 1458 -347
rect 1564 -381 1576 -347
rect 1682 -381 1694 -347
rect 1800 -381 1812 -347
rect 1918 -381 1930 -347
rect 2036 -381 2048 -347
rect 2154 -381 2166 -347
rect 2272 -381 2284 -347
rect 2390 -381 2402 -347
rect 2508 -381 2520 -347
rect 2626 -381 2638 -347
rect 2744 -381 2756 -347
rect 2862 -381 2874 -347
rect -2920 -387 -2862 -381
rect -2802 -387 -2744 -381
rect -2684 -387 -2626 -381
rect -2566 -387 -2508 -381
rect -2448 -387 -2390 -381
rect -2330 -387 -2272 -381
rect -2212 -387 -2154 -381
rect -2094 -387 -2036 -381
rect -1976 -387 -1918 -381
rect -1858 -387 -1800 -381
rect -1740 -387 -1682 -381
rect -1622 -387 -1564 -381
rect -1504 -387 -1446 -381
rect -1386 -387 -1328 -381
rect -1268 -387 -1210 -381
rect -1150 -387 -1092 -381
rect -1032 -387 -974 -381
rect -914 -387 -856 -381
rect -796 -387 -738 -381
rect -678 -387 -620 -381
rect -560 -387 -502 -381
rect -442 -387 -384 -381
rect -324 -387 -266 -381
rect -206 -387 -148 -381
rect -88 -387 -30 -381
rect 30 -387 88 -381
rect 148 -387 206 -381
rect 266 -387 324 -381
rect 384 -387 442 -381
rect 502 -387 560 -381
rect 620 -387 678 -381
rect 738 -387 796 -381
rect 856 -387 914 -381
rect 974 -387 1032 -381
rect 1092 -387 1150 -381
rect 1210 -387 1268 -381
rect 1328 -387 1386 -381
rect 1446 -387 1504 -381
rect 1564 -387 1622 -381
rect 1682 -387 1740 -381
rect 1800 -387 1858 -381
rect 1918 -387 1976 -381
rect 2036 -387 2094 -381
rect 2154 -387 2212 -381
rect 2272 -387 2330 -381
rect 2390 -387 2448 -381
rect 2508 -387 2566 -381
rect 2626 -387 2684 -381
rect 2744 -387 2802 -381
rect 2862 -387 2920 -381
rect -2920 -455 -2862 -449
rect -2802 -455 -2744 -449
rect -2684 -455 -2626 -449
rect -2566 -455 -2508 -449
rect -2448 -455 -2390 -449
rect -2330 -455 -2272 -449
rect -2212 -455 -2154 -449
rect -2094 -455 -2036 -449
rect -1976 -455 -1918 -449
rect -1858 -455 -1800 -449
rect -1740 -455 -1682 -449
rect -1622 -455 -1564 -449
rect -1504 -455 -1446 -449
rect -1386 -455 -1328 -449
rect -1268 -455 -1210 -449
rect -1150 -455 -1092 -449
rect -1032 -455 -974 -449
rect -914 -455 -856 -449
rect -796 -455 -738 -449
rect -678 -455 -620 -449
rect -560 -455 -502 -449
rect -442 -455 -384 -449
rect -324 -455 -266 -449
rect -206 -455 -148 -449
rect -88 -455 -30 -449
rect 30 -455 88 -449
rect 148 -455 206 -449
rect 266 -455 324 -449
rect 384 -455 442 -449
rect 502 -455 560 -449
rect 620 -455 678 -449
rect 738 -455 796 -449
rect 856 -455 914 -449
rect 974 -455 1032 -449
rect 1092 -455 1150 -449
rect 1210 -455 1268 -449
rect 1328 -455 1386 -449
rect 1446 -455 1504 -449
rect 1564 -455 1622 -449
rect 1682 -455 1740 -449
rect 1800 -455 1858 -449
rect 1918 -455 1976 -449
rect 2036 -455 2094 -449
rect 2154 -455 2212 -449
rect 2272 -455 2330 -449
rect 2390 -455 2448 -449
rect 2508 -455 2566 -449
rect 2626 -455 2684 -449
rect 2744 -455 2802 -449
rect 2862 -455 2920 -449
rect -2920 -489 -2908 -455
rect -2802 -489 -2790 -455
rect -2684 -489 -2672 -455
rect -2566 -489 -2554 -455
rect -2448 -489 -2436 -455
rect -2330 -489 -2318 -455
rect -2212 -489 -2200 -455
rect -2094 -489 -2082 -455
rect -1976 -489 -1964 -455
rect -1858 -489 -1846 -455
rect -1740 -489 -1728 -455
rect -1622 -489 -1610 -455
rect -1504 -489 -1492 -455
rect -1386 -489 -1374 -455
rect -1268 -489 -1256 -455
rect -1150 -489 -1138 -455
rect -1032 -489 -1020 -455
rect -914 -489 -902 -455
rect -796 -489 -784 -455
rect -678 -489 -666 -455
rect -560 -489 -548 -455
rect -442 -489 -430 -455
rect -324 -489 -312 -455
rect -206 -489 -194 -455
rect -88 -489 -76 -455
rect 30 -489 42 -455
rect 148 -489 160 -455
rect 266 -489 278 -455
rect 384 -489 396 -455
rect 502 -489 514 -455
rect 620 -489 632 -455
rect 738 -489 750 -455
rect 856 -489 868 -455
rect 974 -489 986 -455
rect 1092 -489 1104 -455
rect 1210 -489 1222 -455
rect 1328 -489 1340 -455
rect 1446 -489 1458 -455
rect 1564 -489 1576 -455
rect 1682 -489 1694 -455
rect 1800 -489 1812 -455
rect 1918 -489 1930 -455
rect 2036 -489 2048 -455
rect 2154 -489 2166 -455
rect 2272 -489 2284 -455
rect 2390 -489 2402 -455
rect 2508 -489 2520 -455
rect 2626 -489 2638 -455
rect 2744 -489 2756 -455
rect 2862 -489 2874 -455
rect -2920 -495 -2862 -489
rect -2802 -495 -2744 -489
rect -2684 -495 -2626 -489
rect -2566 -495 -2508 -489
rect -2448 -495 -2390 -489
rect -2330 -495 -2272 -489
rect -2212 -495 -2154 -489
rect -2094 -495 -2036 -489
rect -1976 -495 -1918 -489
rect -1858 -495 -1800 -489
rect -1740 -495 -1682 -489
rect -1622 -495 -1564 -489
rect -1504 -495 -1446 -489
rect -1386 -495 -1328 -489
rect -1268 -495 -1210 -489
rect -1150 -495 -1092 -489
rect -1032 -495 -974 -489
rect -914 -495 -856 -489
rect -796 -495 -738 -489
rect -678 -495 -620 -489
rect -560 -495 -502 -489
rect -442 -495 -384 -489
rect -324 -495 -266 -489
rect -206 -495 -148 -489
rect -88 -495 -30 -489
rect 30 -495 88 -489
rect 148 -495 206 -489
rect 266 -495 324 -489
rect 384 -495 442 -489
rect 502 -495 560 -489
rect 620 -495 678 -489
rect 738 -495 796 -489
rect 856 -495 914 -489
rect 974 -495 1032 -489
rect 1092 -495 1150 -489
rect 1210 -495 1268 -489
rect 1328 -495 1386 -489
rect 1446 -495 1504 -489
rect 1564 -495 1622 -489
rect 1682 -495 1740 -489
rect 1800 -495 1858 -489
rect 1918 -495 1976 -489
rect 2036 -495 2094 -489
rect 2154 -495 2212 -489
rect 2272 -495 2330 -489
rect 2390 -495 2448 -489
rect 2508 -495 2566 -489
rect 2626 -495 2684 -489
rect 2744 -495 2802 -489
rect 2862 -495 2920 -489
rect -2920 -1183 -2862 -1177
rect -2802 -1183 -2744 -1177
rect -2684 -1183 -2626 -1177
rect -2566 -1183 -2508 -1177
rect -2448 -1183 -2390 -1177
rect -2330 -1183 -2272 -1177
rect -2212 -1183 -2154 -1177
rect -2094 -1183 -2036 -1177
rect -1976 -1183 -1918 -1177
rect -1858 -1183 -1800 -1177
rect -1740 -1183 -1682 -1177
rect -1622 -1183 -1564 -1177
rect -1504 -1183 -1446 -1177
rect -1386 -1183 -1328 -1177
rect -1268 -1183 -1210 -1177
rect -1150 -1183 -1092 -1177
rect -1032 -1183 -974 -1177
rect -914 -1183 -856 -1177
rect -796 -1183 -738 -1177
rect -678 -1183 -620 -1177
rect -560 -1183 -502 -1177
rect -442 -1183 -384 -1177
rect -324 -1183 -266 -1177
rect -206 -1183 -148 -1177
rect -88 -1183 -30 -1177
rect 30 -1183 88 -1177
rect 148 -1183 206 -1177
rect 266 -1183 324 -1177
rect 384 -1183 442 -1177
rect 502 -1183 560 -1177
rect 620 -1183 678 -1177
rect 738 -1183 796 -1177
rect 856 -1183 914 -1177
rect 974 -1183 1032 -1177
rect 1092 -1183 1150 -1177
rect 1210 -1183 1268 -1177
rect 1328 -1183 1386 -1177
rect 1446 -1183 1504 -1177
rect 1564 -1183 1622 -1177
rect 1682 -1183 1740 -1177
rect 1800 -1183 1858 -1177
rect 1918 -1183 1976 -1177
rect 2036 -1183 2094 -1177
rect 2154 -1183 2212 -1177
rect 2272 -1183 2330 -1177
rect 2390 -1183 2448 -1177
rect 2508 -1183 2566 -1177
rect 2626 -1183 2684 -1177
rect 2744 -1183 2802 -1177
rect 2862 -1183 2920 -1177
rect -2920 -1217 -2908 -1183
rect -2802 -1217 -2790 -1183
rect -2684 -1217 -2672 -1183
rect -2566 -1217 -2554 -1183
rect -2448 -1217 -2436 -1183
rect -2330 -1217 -2318 -1183
rect -2212 -1217 -2200 -1183
rect -2094 -1217 -2082 -1183
rect -1976 -1217 -1964 -1183
rect -1858 -1217 -1846 -1183
rect -1740 -1217 -1728 -1183
rect -1622 -1217 -1610 -1183
rect -1504 -1217 -1492 -1183
rect -1386 -1217 -1374 -1183
rect -1268 -1217 -1256 -1183
rect -1150 -1217 -1138 -1183
rect -1032 -1217 -1020 -1183
rect -914 -1217 -902 -1183
rect -796 -1217 -784 -1183
rect -678 -1217 -666 -1183
rect -560 -1217 -548 -1183
rect -442 -1217 -430 -1183
rect -324 -1217 -312 -1183
rect -206 -1217 -194 -1183
rect -88 -1217 -76 -1183
rect 30 -1217 42 -1183
rect 148 -1217 160 -1183
rect 266 -1217 278 -1183
rect 384 -1217 396 -1183
rect 502 -1217 514 -1183
rect 620 -1217 632 -1183
rect 738 -1217 750 -1183
rect 856 -1217 868 -1183
rect 974 -1217 986 -1183
rect 1092 -1217 1104 -1183
rect 1210 -1217 1222 -1183
rect 1328 -1217 1340 -1183
rect 1446 -1217 1458 -1183
rect 1564 -1217 1576 -1183
rect 1682 -1217 1694 -1183
rect 1800 -1217 1812 -1183
rect 1918 -1217 1930 -1183
rect 2036 -1217 2048 -1183
rect 2154 -1217 2166 -1183
rect 2272 -1217 2284 -1183
rect 2390 -1217 2402 -1183
rect 2508 -1217 2520 -1183
rect 2626 -1217 2638 -1183
rect 2744 -1217 2756 -1183
rect 2862 -1217 2874 -1183
rect -2920 -1223 -2862 -1217
rect -2802 -1223 -2744 -1217
rect -2684 -1223 -2626 -1217
rect -2566 -1223 -2508 -1217
rect -2448 -1223 -2390 -1217
rect -2330 -1223 -2272 -1217
rect -2212 -1223 -2154 -1217
rect -2094 -1223 -2036 -1217
rect -1976 -1223 -1918 -1217
rect -1858 -1223 -1800 -1217
rect -1740 -1223 -1682 -1217
rect -1622 -1223 -1564 -1217
rect -1504 -1223 -1446 -1217
rect -1386 -1223 -1328 -1217
rect -1268 -1223 -1210 -1217
rect -1150 -1223 -1092 -1217
rect -1032 -1223 -974 -1217
rect -914 -1223 -856 -1217
rect -796 -1223 -738 -1217
rect -678 -1223 -620 -1217
rect -560 -1223 -502 -1217
rect -442 -1223 -384 -1217
rect -324 -1223 -266 -1217
rect -206 -1223 -148 -1217
rect -88 -1223 -30 -1217
rect 30 -1223 88 -1217
rect 148 -1223 206 -1217
rect 266 -1223 324 -1217
rect 384 -1223 442 -1217
rect 502 -1223 560 -1217
rect 620 -1223 678 -1217
rect 738 -1223 796 -1217
rect 856 -1223 914 -1217
rect 974 -1223 1032 -1217
rect 1092 -1223 1150 -1217
rect 1210 -1223 1268 -1217
rect 1328 -1223 1386 -1217
rect 1446 -1223 1504 -1217
rect 1564 -1223 1622 -1217
rect 1682 -1223 1740 -1217
rect 1800 -1223 1858 -1217
rect 1918 -1223 1976 -1217
rect 2036 -1223 2094 -1217
rect 2154 -1223 2212 -1217
rect 2272 -1223 2330 -1217
rect 2390 -1223 2448 -1217
rect 2508 -1223 2566 -1217
rect 2626 -1223 2684 -1217
rect 2744 -1223 2802 -1217
rect 2862 -1223 2920 -1217
<< nwell >>
rect -3117 -1355 3117 1355
<< pmos >>
rect -2921 536 -2861 1136
rect -2803 536 -2743 1136
rect -2685 536 -2625 1136
rect -2567 536 -2507 1136
rect -2449 536 -2389 1136
rect -2331 536 -2271 1136
rect -2213 536 -2153 1136
rect -2095 536 -2035 1136
rect -1977 536 -1917 1136
rect -1859 536 -1799 1136
rect -1741 536 -1681 1136
rect -1623 536 -1563 1136
rect -1505 536 -1445 1136
rect -1387 536 -1327 1136
rect -1269 536 -1209 1136
rect -1151 536 -1091 1136
rect -1033 536 -973 1136
rect -915 536 -855 1136
rect -797 536 -737 1136
rect -679 536 -619 1136
rect -561 536 -501 1136
rect -443 536 -383 1136
rect -325 536 -265 1136
rect -207 536 -147 1136
rect -89 536 -29 1136
rect 29 536 89 1136
rect 147 536 207 1136
rect 265 536 325 1136
rect 383 536 443 1136
rect 501 536 561 1136
rect 619 536 679 1136
rect 737 536 797 1136
rect 855 536 915 1136
rect 973 536 1033 1136
rect 1091 536 1151 1136
rect 1209 536 1269 1136
rect 1327 536 1387 1136
rect 1445 536 1505 1136
rect 1563 536 1623 1136
rect 1681 536 1741 1136
rect 1799 536 1859 1136
rect 1917 536 1977 1136
rect 2035 536 2095 1136
rect 2153 536 2213 1136
rect 2271 536 2331 1136
rect 2389 536 2449 1136
rect 2507 536 2567 1136
rect 2625 536 2685 1136
rect 2743 536 2803 1136
rect 2861 536 2921 1136
rect -2921 -300 -2861 300
rect -2803 -300 -2743 300
rect -2685 -300 -2625 300
rect -2567 -300 -2507 300
rect -2449 -300 -2389 300
rect -2331 -300 -2271 300
rect -2213 -300 -2153 300
rect -2095 -300 -2035 300
rect -1977 -300 -1917 300
rect -1859 -300 -1799 300
rect -1741 -300 -1681 300
rect -1623 -300 -1563 300
rect -1505 -300 -1445 300
rect -1387 -300 -1327 300
rect -1269 -300 -1209 300
rect -1151 -300 -1091 300
rect -1033 -300 -973 300
rect -915 -300 -855 300
rect -797 -300 -737 300
rect -679 -300 -619 300
rect -561 -300 -501 300
rect -443 -300 -383 300
rect -325 -300 -265 300
rect -207 -300 -147 300
rect -89 -300 -29 300
rect 29 -300 89 300
rect 147 -300 207 300
rect 265 -300 325 300
rect 383 -300 443 300
rect 501 -300 561 300
rect 619 -300 679 300
rect 737 -300 797 300
rect 855 -300 915 300
rect 973 -300 1033 300
rect 1091 -300 1151 300
rect 1209 -300 1269 300
rect 1327 -300 1387 300
rect 1445 -300 1505 300
rect 1563 -300 1623 300
rect 1681 -300 1741 300
rect 1799 -300 1859 300
rect 1917 -300 1977 300
rect 2035 -300 2095 300
rect 2153 -300 2213 300
rect 2271 -300 2331 300
rect 2389 -300 2449 300
rect 2507 -300 2567 300
rect 2625 -300 2685 300
rect 2743 -300 2803 300
rect 2861 -300 2921 300
rect -2921 -1136 -2861 -536
rect -2803 -1136 -2743 -536
rect -2685 -1136 -2625 -536
rect -2567 -1136 -2507 -536
rect -2449 -1136 -2389 -536
rect -2331 -1136 -2271 -536
rect -2213 -1136 -2153 -536
rect -2095 -1136 -2035 -536
rect -1977 -1136 -1917 -536
rect -1859 -1136 -1799 -536
rect -1741 -1136 -1681 -536
rect -1623 -1136 -1563 -536
rect -1505 -1136 -1445 -536
rect -1387 -1136 -1327 -536
rect -1269 -1136 -1209 -536
rect -1151 -1136 -1091 -536
rect -1033 -1136 -973 -536
rect -915 -1136 -855 -536
rect -797 -1136 -737 -536
rect -679 -1136 -619 -536
rect -561 -1136 -501 -536
rect -443 -1136 -383 -536
rect -325 -1136 -265 -536
rect -207 -1136 -147 -536
rect -89 -1136 -29 -536
rect 29 -1136 89 -536
rect 147 -1136 207 -536
rect 265 -1136 325 -536
rect 383 -1136 443 -536
rect 501 -1136 561 -536
rect 619 -1136 679 -536
rect 737 -1136 797 -536
rect 855 -1136 915 -536
rect 973 -1136 1033 -536
rect 1091 -1136 1151 -536
rect 1209 -1136 1269 -536
rect 1327 -1136 1387 -536
rect 1445 -1136 1505 -536
rect 1563 -1136 1623 -536
rect 1681 -1136 1741 -536
rect 1799 -1136 1859 -536
rect 1917 -1136 1977 -536
rect 2035 -1136 2095 -536
rect 2153 -1136 2213 -536
rect 2271 -1136 2331 -536
rect 2389 -1136 2449 -536
rect 2507 -1136 2567 -536
rect 2625 -1136 2685 -536
rect 2743 -1136 2803 -536
rect 2861 -1136 2921 -536
<< pdiff >>
rect -2979 1124 -2921 1136
rect -2979 548 -2967 1124
rect -2933 548 -2921 1124
rect -2979 536 -2921 548
rect -2861 1124 -2803 1136
rect -2861 548 -2849 1124
rect -2815 548 -2803 1124
rect -2861 536 -2803 548
rect -2743 1124 -2685 1136
rect -2743 548 -2731 1124
rect -2697 548 -2685 1124
rect -2743 536 -2685 548
rect -2625 1124 -2567 1136
rect -2625 548 -2613 1124
rect -2579 548 -2567 1124
rect -2625 536 -2567 548
rect -2507 1124 -2449 1136
rect -2507 548 -2495 1124
rect -2461 548 -2449 1124
rect -2507 536 -2449 548
rect -2389 1124 -2331 1136
rect -2389 548 -2377 1124
rect -2343 548 -2331 1124
rect -2389 536 -2331 548
rect -2271 1124 -2213 1136
rect -2271 548 -2259 1124
rect -2225 548 -2213 1124
rect -2271 536 -2213 548
rect -2153 1124 -2095 1136
rect -2153 548 -2141 1124
rect -2107 548 -2095 1124
rect -2153 536 -2095 548
rect -2035 1124 -1977 1136
rect -2035 548 -2023 1124
rect -1989 548 -1977 1124
rect -2035 536 -1977 548
rect -1917 1124 -1859 1136
rect -1917 548 -1905 1124
rect -1871 548 -1859 1124
rect -1917 536 -1859 548
rect -1799 1124 -1741 1136
rect -1799 548 -1787 1124
rect -1753 548 -1741 1124
rect -1799 536 -1741 548
rect -1681 1124 -1623 1136
rect -1681 548 -1669 1124
rect -1635 548 -1623 1124
rect -1681 536 -1623 548
rect -1563 1124 -1505 1136
rect -1563 548 -1551 1124
rect -1517 548 -1505 1124
rect -1563 536 -1505 548
rect -1445 1124 -1387 1136
rect -1445 548 -1433 1124
rect -1399 548 -1387 1124
rect -1445 536 -1387 548
rect -1327 1124 -1269 1136
rect -1327 548 -1315 1124
rect -1281 548 -1269 1124
rect -1327 536 -1269 548
rect -1209 1124 -1151 1136
rect -1209 548 -1197 1124
rect -1163 548 -1151 1124
rect -1209 536 -1151 548
rect -1091 1124 -1033 1136
rect -1091 548 -1079 1124
rect -1045 548 -1033 1124
rect -1091 536 -1033 548
rect -973 1124 -915 1136
rect -973 548 -961 1124
rect -927 548 -915 1124
rect -973 536 -915 548
rect -855 1124 -797 1136
rect -855 548 -843 1124
rect -809 548 -797 1124
rect -855 536 -797 548
rect -737 1124 -679 1136
rect -737 548 -725 1124
rect -691 548 -679 1124
rect -737 536 -679 548
rect -619 1124 -561 1136
rect -619 548 -607 1124
rect -573 548 -561 1124
rect -619 536 -561 548
rect -501 1124 -443 1136
rect -501 548 -489 1124
rect -455 548 -443 1124
rect -501 536 -443 548
rect -383 1124 -325 1136
rect -383 548 -371 1124
rect -337 548 -325 1124
rect -383 536 -325 548
rect -265 1124 -207 1136
rect -265 548 -253 1124
rect -219 548 -207 1124
rect -265 536 -207 548
rect -147 1124 -89 1136
rect -147 548 -135 1124
rect -101 548 -89 1124
rect -147 536 -89 548
rect -29 1124 29 1136
rect -29 548 -17 1124
rect 17 548 29 1124
rect -29 536 29 548
rect 89 1124 147 1136
rect 89 548 101 1124
rect 135 548 147 1124
rect 89 536 147 548
rect 207 1124 265 1136
rect 207 548 219 1124
rect 253 548 265 1124
rect 207 536 265 548
rect 325 1124 383 1136
rect 325 548 337 1124
rect 371 548 383 1124
rect 325 536 383 548
rect 443 1124 501 1136
rect 443 548 455 1124
rect 489 548 501 1124
rect 443 536 501 548
rect 561 1124 619 1136
rect 561 548 573 1124
rect 607 548 619 1124
rect 561 536 619 548
rect 679 1124 737 1136
rect 679 548 691 1124
rect 725 548 737 1124
rect 679 536 737 548
rect 797 1124 855 1136
rect 797 548 809 1124
rect 843 548 855 1124
rect 797 536 855 548
rect 915 1124 973 1136
rect 915 548 927 1124
rect 961 548 973 1124
rect 915 536 973 548
rect 1033 1124 1091 1136
rect 1033 548 1045 1124
rect 1079 548 1091 1124
rect 1033 536 1091 548
rect 1151 1124 1209 1136
rect 1151 548 1163 1124
rect 1197 548 1209 1124
rect 1151 536 1209 548
rect 1269 1124 1327 1136
rect 1269 548 1281 1124
rect 1315 548 1327 1124
rect 1269 536 1327 548
rect 1387 1124 1445 1136
rect 1387 548 1399 1124
rect 1433 548 1445 1124
rect 1387 536 1445 548
rect 1505 1124 1563 1136
rect 1505 548 1517 1124
rect 1551 548 1563 1124
rect 1505 536 1563 548
rect 1623 1124 1681 1136
rect 1623 548 1635 1124
rect 1669 548 1681 1124
rect 1623 536 1681 548
rect 1741 1124 1799 1136
rect 1741 548 1753 1124
rect 1787 548 1799 1124
rect 1741 536 1799 548
rect 1859 1124 1917 1136
rect 1859 548 1871 1124
rect 1905 548 1917 1124
rect 1859 536 1917 548
rect 1977 1124 2035 1136
rect 1977 548 1989 1124
rect 2023 548 2035 1124
rect 1977 536 2035 548
rect 2095 1124 2153 1136
rect 2095 548 2107 1124
rect 2141 548 2153 1124
rect 2095 536 2153 548
rect 2213 1124 2271 1136
rect 2213 548 2225 1124
rect 2259 548 2271 1124
rect 2213 536 2271 548
rect 2331 1124 2389 1136
rect 2331 548 2343 1124
rect 2377 548 2389 1124
rect 2331 536 2389 548
rect 2449 1124 2507 1136
rect 2449 548 2461 1124
rect 2495 548 2507 1124
rect 2449 536 2507 548
rect 2567 1124 2625 1136
rect 2567 548 2579 1124
rect 2613 548 2625 1124
rect 2567 536 2625 548
rect 2685 1124 2743 1136
rect 2685 548 2697 1124
rect 2731 548 2743 1124
rect 2685 536 2743 548
rect 2803 1124 2861 1136
rect 2803 548 2815 1124
rect 2849 548 2861 1124
rect 2803 536 2861 548
rect 2921 1124 2979 1136
rect 2921 548 2933 1124
rect 2967 548 2979 1124
rect 2921 536 2979 548
rect -2979 288 -2921 300
rect -2979 -288 -2967 288
rect -2933 -288 -2921 288
rect -2979 -300 -2921 -288
rect -2861 288 -2803 300
rect -2861 -288 -2849 288
rect -2815 -288 -2803 288
rect -2861 -300 -2803 -288
rect -2743 288 -2685 300
rect -2743 -288 -2731 288
rect -2697 -288 -2685 288
rect -2743 -300 -2685 -288
rect -2625 288 -2567 300
rect -2625 -288 -2613 288
rect -2579 -288 -2567 288
rect -2625 -300 -2567 -288
rect -2507 288 -2449 300
rect -2507 -288 -2495 288
rect -2461 -288 -2449 288
rect -2507 -300 -2449 -288
rect -2389 288 -2331 300
rect -2389 -288 -2377 288
rect -2343 -288 -2331 288
rect -2389 -300 -2331 -288
rect -2271 288 -2213 300
rect -2271 -288 -2259 288
rect -2225 -288 -2213 288
rect -2271 -300 -2213 -288
rect -2153 288 -2095 300
rect -2153 -288 -2141 288
rect -2107 -288 -2095 288
rect -2153 -300 -2095 -288
rect -2035 288 -1977 300
rect -2035 -288 -2023 288
rect -1989 -288 -1977 288
rect -2035 -300 -1977 -288
rect -1917 288 -1859 300
rect -1917 -288 -1905 288
rect -1871 -288 -1859 288
rect -1917 -300 -1859 -288
rect -1799 288 -1741 300
rect -1799 -288 -1787 288
rect -1753 -288 -1741 288
rect -1799 -300 -1741 -288
rect -1681 288 -1623 300
rect -1681 -288 -1669 288
rect -1635 -288 -1623 288
rect -1681 -300 -1623 -288
rect -1563 288 -1505 300
rect -1563 -288 -1551 288
rect -1517 -288 -1505 288
rect -1563 -300 -1505 -288
rect -1445 288 -1387 300
rect -1445 -288 -1433 288
rect -1399 -288 -1387 288
rect -1445 -300 -1387 -288
rect -1327 288 -1269 300
rect -1327 -288 -1315 288
rect -1281 -288 -1269 288
rect -1327 -300 -1269 -288
rect -1209 288 -1151 300
rect -1209 -288 -1197 288
rect -1163 -288 -1151 288
rect -1209 -300 -1151 -288
rect -1091 288 -1033 300
rect -1091 -288 -1079 288
rect -1045 -288 -1033 288
rect -1091 -300 -1033 -288
rect -973 288 -915 300
rect -973 -288 -961 288
rect -927 -288 -915 288
rect -973 -300 -915 -288
rect -855 288 -797 300
rect -855 -288 -843 288
rect -809 -288 -797 288
rect -855 -300 -797 -288
rect -737 288 -679 300
rect -737 -288 -725 288
rect -691 -288 -679 288
rect -737 -300 -679 -288
rect -619 288 -561 300
rect -619 -288 -607 288
rect -573 -288 -561 288
rect -619 -300 -561 -288
rect -501 288 -443 300
rect -501 -288 -489 288
rect -455 -288 -443 288
rect -501 -300 -443 -288
rect -383 288 -325 300
rect -383 -288 -371 288
rect -337 -288 -325 288
rect -383 -300 -325 -288
rect -265 288 -207 300
rect -265 -288 -253 288
rect -219 -288 -207 288
rect -265 -300 -207 -288
rect -147 288 -89 300
rect -147 -288 -135 288
rect -101 -288 -89 288
rect -147 -300 -89 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 89 288 147 300
rect 89 -288 101 288
rect 135 -288 147 288
rect 89 -300 147 -288
rect 207 288 265 300
rect 207 -288 219 288
rect 253 -288 265 288
rect 207 -300 265 -288
rect 325 288 383 300
rect 325 -288 337 288
rect 371 -288 383 288
rect 325 -300 383 -288
rect 443 288 501 300
rect 443 -288 455 288
rect 489 -288 501 288
rect 443 -300 501 -288
rect 561 288 619 300
rect 561 -288 573 288
rect 607 -288 619 288
rect 561 -300 619 -288
rect 679 288 737 300
rect 679 -288 691 288
rect 725 -288 737 288
rect 679 -300 737 -288
rect 797 288 855 300
rect 797 -288 809 288
rect 843 -288 855 288
rect 797 -300 855 -288
rect 915 288 973 300
rect 915 -288 927 288
rect 961 -288 973 288
rect 915 -300 973 -288
rect 1033 288 1091 300
rect 1033 -288 1045 288
rect 1079 -288 1091 288
rect 1033 -300 1091 -288
rect 1151 288 1209 300
rect 1151 -288 1163 288
rect 1197 -288 1209 288
rect 1151 -300 1209 -288
rect 1269 288 1327 300
rect 1269 -288 1281 288
rect 1315 -288 1327 288
rect 1269 -300 1327 -288
rect 1387 288 1445 300
rect 1387 -288 1399 288
rect 1433 -288 1445 288
rect 1387 -300 1445 -288
rect 1505 288 1563 300
rect 1505 -288 1517 288
rect 1551 -288 1563 288
rect 1505 -300 1563 -288
rect 1623 288 1681 300
rect 1623 -288 1635 288
rect 1669 -288 1681 288
rect 1623 -300 1681 -288
rect 1741 288 1799 300
rect 1741 -288 1753 288
rect 1787 -288 1799 288
rect 1741 -300 1799 -288
rect 1859 288 1917 300
rect 1859 -288 1871 288
rect 1905 -288 1917 288
rect 1859 -300 1917 -288
rect 1977 288 2035 300
rect 1977 -288 1989 288
rect 2023 -288 2035 288
rect 1977 -300 2035 -288
rect 2095 288 2153 300
rect 2095 -288 2107 288
rect 2141 -288 2153 288
rect 2095 -300 2153 -288
rect 2213 288 2271 300
rect 2213 -288 2225 288
rect 2259 -288 2271 288
rect 2213 -300 2271 -288
rect 2331 288 2389 300
rect 2331 -288 2343 288
rect 2377 -288 2389 288
rect 2331 -300 2389 -288
rect 2449 288 2507 300
rect 2449 -288 2461 288
rect 2495 -288 2507 288
rect 2449 -300 2507 -288
rect 2567 288 2625 300
rect 2567 -288 2579 288
rect 2613 -288 2625 288
rect 2567 -300 2625 -288
rect 2685 288 2743 300
rect 2685 -288 2697 288
rect 2731 -288 2743 288
rect 2685 -300 2743 -288
rect 2803 288 2861 300
rect 2803 -288 2815 288
rect 2849 -288 2861 288
rect 2803 -300 2861 -288
rect 2921 288 2979 300
rect 2921 -288 2933 288
rect 2967 -288 2979 288
rect 2921 -300 2979 -288
rect -2979 -548 -2921 -536
rect -2979 -1124 -2967 -548
rect -2933 -1124 -2921 -548
rect -2979 -1136 -2921 -1124
rect -2861 -548 -2803 -536
rect -2861 -1124 -2849 -548
rect -2815 -1124 -2803 -548
rect -2861 -1136 -2803 -1124
rect -2743 -548 -2685 -536
rect -2743 -1124 -2731 -548
rect -2697 -1124 -2685 -548
rect -2743 -1136 -2685 -1124
rect -2625 -548 -2567 -536
rect -2625 -1124 -2613 -548
rect -2579 -1124 -2567 -548
rect -2625 -1136 -2567 -1124
rect -2507 -548 -2449 -536
rect -2507 -1124 -2495 -548
rect -2461 -1124 -2449 -548
rect -2507 -1136 -2449 -1124
rect -2389 -548 -2331 -536
rect -2389 -1124 -2377 -548
rect -2343 -1124 -2331 -548
rect -2389 -1136 -2331 -1124
rect -2271 -548 -2213 -536
rect -2271 -1124 -2259 -548
rect -2225 -1124 -2213 -548
rect -2271 -1136 -2213 -1124
rect -2153 -548 -2095 -536
rect -2153 -1124 -2141 -548
rect -2107 -1124 -2095 -548
rect -2153 -1136 -2095 -1124
rect -2035 -548 -1977 -536
rect -2035 -1124 -2023 -548
rect -1989 -1124 -1977 -548
rect -2035 -1136 -1977 -1124
rect -1917 -548 -1859 -536
rect -1917 -1124 -1905 -548
rect -1871 -1124 -1859 -548
rect -1917 -1136 -1859 -1124
rect -1799 -548 -1741 -536
rect -1799 -1124 -1787 -548
rect -1753 -1124 -1741 -548
rect -1799 -1136 -1741 -1124
rect -1681 -548 -1623 -536
rect -1681 -1124 -1669 -548
rect -1635 -1124 -1623 -548
rect -1681 -1136 -1623 -1124
rect -1563 -548 -1505 -536
rect -1563 -1124 -1551 -548
rect -1517 -1124 -1505 -548
rect -1563 -1136 -1505 -1124
rect -1445 -548 -1387 -536
rect -1445 -1124 -1433 -548
rect -1399 -1124 -1387 -548
rect -1445 -1136 -1387 -1124
rect -1327 -548 -1269 -536
rect -1327 -1124 -1315 -548
rect -1281 -1124 -1269 -548
rect -1327 -1136 -1269 -1124
rect -1209 -548 -1151 -536
rect -1209 -1124 -1197 -548
rect -1163 -1124 -1151 -548
rect -1209 -1136 -1151 -1124
rect -1091 -548 -1033 -536
rect -1091 -1124 -1079 -548
rect -1045 -1124 -1033 -548
rect -1091 -1136 -1033 -1124
rect -973 -548 -915 -536
rect -973 -1124 -961 -548
rect -927 -1124 -915 -548
rect -973 -1136 -915 -1124
rect -855 -548 -797 -536
rect -855 -1124 -843 -548
rect -809 -1124 -797 -548
rect -855 -1136 -797 -1124
rect -737 -548 -679 -536
rect -737 -1124 -725 -548
rect -691 -1124 -679 -548
rect -737 -1136 -679 -1124
rect -619 -548 -561 -536
rect -619 -1124 -607 -548
rect -573 -1124 -561 -548
rect -619 -1136 -561 -1124
rect -501 -548 -443 -536
rect -501 -1124 -489 -548
rect -455 -1124 -443 -548
rect -501 -1136 -443 -1124
rect -383 -548 -325 -536
rect -383 -1124 -371 -548
rect -337 -1124 -325 -548
rect -383 -1136 -325 -1124
rect -265 -548 -207 -536
rect -265 -1124 -253 -548
rect -219 -1124 -207 -548
rect -265 -1136 -207 -1124
rect -147 -548 -89 -536
rect -147 -1124 -135 -548
rect -101 -1124 -89 -548
rect -147 -1136 -89 -1124
rect -29 -548 29 -536
rect -29 -1124 -17 -548
rect 17 -1124 29 -548
rect -29 -1136 29 -1124
rect 89 -548 147 -536
rect 89 -1124 101 -548
rect 135 -1124 147 -548
rect 89 -1136 147 -1124
rect 207 -548 265 -536
rect 207 -1124 219 -548
rect 253 -1124 265 -548
rect 207 -1136 265 -1124
rect 325 -548 383 -536
rect 325 -1124 337 -548
rect 371 -1124 383 -548
rect 325 -1136 383 -1124
rect 443 -548 501 -536
rect 443 -1124 455 -548
rect 489 -1124 501 -548
rect 443 -1136 501 -1124
rect 561 -548 619 -536
rect 561 -1124 573 -548
rect 607 -1124 619 -548
rect 561 -1136 619 -1124
rect 679 -548 737 -536
rect 679 -1124 691 -548
rect 725 -1124 737 -548
rect 679 -1136 737 -1124
rect 797 -548 855 -536
rect 797 -1124 809 -548
rect 843 -1124 855 -548
rect 797 -1136 855 -1124
rect 915 -548 973 -536
rect 915 -1124 927 -548
rect 961 -1124 973 -548
rect 915 -1136 973 -1124
rect 1033 -548 1091 -536
rect 1033 -1124 1045 -548
rect 1079 -1124 1091 -548
rect 1033 -1136 1091 -1124
rect 1151 -548 1209 -536
rect 1151 -1124 1163 -548
rect 1197 -1124 1209 -548
rect 1151 -1136 1209 -1124
rect 1269 -548 1327 -536
rect 1269 -1124 1281 -548
rect 1315 -1124 1327 -548
rect 1269 -1136 1327 -1124
rect 1387 -548 1445 -536
rect 1387 -1124 1399 -548
rect 1433 -1124 1445 -548
rect 1387 -1136 1445 -1124
rect 1505 -548 1563 -536
rect 1505 -1124 1517 -548
rect 1551 -1124 1563 -548
rect 1505 -1136 1563 -1124
rect 1623 -548 1681 -536
rect 1623 -1124 1635 -548
rect 1669 -1124 1681 -548
rect 1623 -1136 1681 -1124
rect 1741 -548 1799 -536
rect 1741 -1124 1753 -548
rect 1787 -1124 1799 -548
rect 1741 -1136 1799 -1124
rect 1859 -548 1917 -536
rect 1859 -1124 1871 -548
rect 1905 -1124 1917 -548
rect 1859 -1136 1917 -1124
rect 1977 -548 2035 -536
rect 1977 -1124 1989 -548
rect 2023 -1124 2035 -548
rect 1977 -1136 2035 -1124
rect 2095 -548 2153 -536
rect 2095 -1124 2107 -548
rect 2141 -1124 2153 -548
rect 2095 -1136 2153 -1124
rect 2213 -548 2271 -536
rect 2213 -1124 2225 -548
rect 2259 -1124 2271 -548
rect 2213 -1136 2271 -1124
rect 2331 -548 2389 -536
rect 2331 -1124 2343 -548
rect 2377 -1124 2389 -548
rect 2331 -1136 2389 -1124
rect 2449 -548 2507 -536
rect 2449 -1124 2461 -548
rect 2495 -1124 2507 -548
rect 2449 -1136 2507 -1124
rect 2567 -548 2625 -536
rect 2567 -1124 2579 -548
rect 2613 -1124 2625 -548
rect 2567 -1136 2625 -1124
rect 2685 -548 2743 -536
rect 2685 -1124 2697 -548
rect 2731 -1124 2743 -548
rect 2685 -1136 2743 -1124
rect 2803 -548 2861 -536
rect 2803 -1124 2815 -548
rect 2849 -1124 2861 -548
rect 2803 -1136 2861 -1124
rect 2921 -548 2979 -536
rect 2921 -1124 2933 -548
rect 2967 -1124 2979 -548
rect 2921 -1136 2979 -1124
<< pdiffc >>
rect -2967 548 -2933 1124
rect -2849 548 -2815 1124
rect -2731 548 -2697 1124
rect -2613 548 -2579 1124
rect -2495 548 -2461 1124
rect -2377 548 -2343 1124
rect -2259 548 -2225 1124
rect -2141 548 -2107 1124
rect -2023 548 -1989 1124
rect -1905 548 -1871 1124
rect -1787 548 -1753 1124
rect -1669 548 -1635 1124
rect -1551 548 -1517 1124
rect -1433 548 -1399 1124
rect -1315 548 -1281 1124
rect -1197 548 -1163 1124
rect -1079 548 -1045 1124
rect -961 548 -927 1124
rect -843 548 -809 1124
rect -725 548 -691 1124
rect -607 548 -573 1124
rect -489 548 -455 1124
rect -371 548 -337 1124
rect -253 548 -219 1124
rect -135 548 -101 1124
rect -17 548 17 1124
rect 101 548 135 1124
rect 219 548 253 1124
rect 337 548 371 1124
rect 455 548 489 1124
rect 573 548 607 1124
rect 691 548 725 1124
rect 809 548 843 1124
rect 927 548 961 1124
rect 1045 548 1079 1124
rect 1163 548 1197 1124
rect 1281 548 1315 1124
rect 1399 548 1433 1124
rect 1517 548 1551 1124
rect 1635 548 1669 1124
rect 1753 548 1787 1124
rect 1871 548 1905 1124
rect 1989 548 2023 1124
rect 2107 548 2141 1124
rect 2225 548 2259 1124
rect 2343 548 2377 1124
rect 2461 548 2495 1124
rect 2579 548 2613 1124
rect 2697 548 2731 1124
rect 2815 548 2849 1124
rect 2933 548 2967 1124
rect -2967 -288 -2933 288
rect -2849 -288 -2815 288
rect -2731 -288 -2697 288
rect -2613 -288 -2579 288
rect -2495 -288 -2461 288
rect -2377 -288 -2343 288
rect -2259 -288 -2225 288
rect -2141 -288 -2107 288
rect -2023 -288 -1989 288
rect -1905 -288 -1871 288
rect -1787 -288 -1753 288
rect -1669 -288 -1635 288
rect -1551 -288 -1517 288
rect -1433 -288 -1399 288
rect -1315 -288 -1281 288
rect -1197 -288 -1163 288
rect -1079 -288 -1045 288
rect -961 -288 -927 288
rect -843 -288 -809 288
rect -725 -288 -691 288
rect -607 -288 -573 288
rect -489 -288 -455 288
rect -371 -288 -337 288
rect -253 -288 -219 288
rect -135 -288 -101 288
rect -17 -288 17 288
rect 101 -288 135 288
rect 219 -288 253 288
rect 337 -288 371 288
rect 455 -288 489 288
rect 573 -288 607 288
rect 691 -288 725 288
rect 809 -288 843 288
rect 927 -288 961 288
rect 1045 -288 1079 288
rect 1163 -288 1197 288
rect 1281 -288 1315 288
rect 1399 -288 1433 288
rect 1517 -288 1551 288
rect 1635 -288 1669 288
rect 1753 -288 1787 288
rect 1871 -288 1905 288
rect 1989 -288 2023 288
rect 2107 -288 2141 288
rect 2225 -288 2259 288
rect 2343 -288 2377 288
rect 2461 -288 2495 288
rect 2579 -288 2613 288
rect 2697 -288 2731 288
rect 2815 -288 2849 288
rect 2933 -288 2967 288
rect -2967 -1124 -2933 -548
rect -2849 -1124 -2815 -548
rect -2731 -1124 -2697 -548
rect -2613 -1124 -2579 -548
rect -2495 -1124 -2461 -548
rect -2377 -1124 -2343 -548
rect -2259 -1124 -2225 -548
rect -2141 -1124 -2107 -548
rect -2023 -1124 -1989 -548
rect -1905 -1124 -1871 -548
rect -1787 -1124 -1753 -548
rect -1669 -1124 -1635 -548
rect -1551 -1124 -1517 -548
rect -1433 -1124 -1399 -548
rect -1315 -1124 -1281 -548
rect -1197 -1124 -1163 -548
rect -1079 -1124 -1045 -548
rect -961 -1124 -927 -548
rect -843 -1124 -809 -548
rect -725 -1124 -691 -548
rect -607 -1124 -573 -548
rect -489 -1124 -455 -548
rect -371 -1124 -337 -548
rect -253 -1124 -219 -548
rect -135 -1124 -101 -548
rect -17 -1124 17 -548
rect 101 -1124 135 -548
rect 219 -1124 253 -548
rect 337 -1124 371 -548
rect 455 -1124 489 -548
rect 573 -1124 607 -548
rect 691 -1124 725 -548
rect 809 -1124 843 -548
rect 927 -1124 961 -548
rect 1045 -1124 1079 -548
rect 1163 -1124 1197 -548
rect 1281 -1124 1315 -548
rect 1399 -1124 1433 -548
rect 1517 -1124 1551 -548
rect 1635 -1124 1669 -548
rect 1753 -1124 1787 -548
rect 1871 -1124 1905 -548
rect 1989 -1124 2023 -548
rect 2107 -1124 2141 -548
rect 2225 -1124 2259 -548
rect 2343 -1124 2377 -548
rect 2461 -1124 2495 -548
rect 2579 -1124 2613 -548
rect 2697 -1124 2731 -548
rect 2815 -1124 2849 -548
rect 2933 -1124 2967 -548
<< nsubdiff >>
rect -3081 1285 -2985 1319
rect 2985 1285 3081 1319
rect -3081 1223 -3047 1285
rect 3047 1223 3081 1285
rect -3081 -1285 -3047 -1223
rect 3047 -1285 3081 -1223
rect -3081 -1319 -2985 -1285
rect 2985 -1319 3081 -1285
<< nsubdiffcont >>
rect -2985 1285 2985 1319
rect -3081 -1223 -3047 1223
rect 3047 -1223 3081 1223
rect -2985 -1319 2985 -1285
<< poly >>
rect -2924 1217 -2858 1233
rect -2924 1183 -2908 1217
rect -2874 1183 -2858 1217
rect -2924 1167 -2858 1183
rect -2806 1217 -2740 1233
rect -2806 1183 -2790 1217
rect -2756 1183 -2740 1217
rect -2806 1167 -2740 1183
rect -2688 1217 -2622 1233
rect -2688 1183 -2672 1217
rect -2638 1183 -2622 1217
rect -2688 1167 -2622 1183
rect -2570 1217 -2504 1233
rect -2570 1183 -2554 1217
rect -2520 1183 -2504 1217
rect -2570 1167 -2504 1183
rect -2452 1217 -2386 1233
rect -2452 1183 -2436 1217
rect -2402 1183 -2386 1217
rect -2452 1167 -2386 1183
rect -2334 1217 -2268 1233
rect -2334 1183 -2318 1217
rect -2284 1183 -2268 1217
rect -2334 1167 -2268 1183
rect -2216 1217 -2150 1233
rect -2216 1183 -2200 1217
rect -2166 1183 -2150 1217
rect -2216 1167 -2150 1183
rect -2098 1217 -2032 1233
rect -2098 1183 -2082 1217
rect -2048 1183 -2032 1217
rect -2098 1167 -2032 1183
rect -1980 1217 -1914 1233
rect -1980 1183 -1964 1217
rect -1930 1183 -1914 1217
rect -1980 1167 -1914 1183
rect -1862 1217 -1796 1233
rect -1862 1183 -1846 1217
rect -1812 1183 -1796 1217
rect -1862 1167 -1796 1183
rect -1744 1217 -1678 1233
rect -1744 1183 -1728 1217
rect -1694 1183 -1678 1217
rect -1744 1167 -1678 1183
rect -1626 1217 -1560 1233
rect -1626 1183 -1610 1217
rect -1576 1183 -1560 1217
rect -1626 1167 -1560 1183
rect -1508 1217 -1442 1233
rect -1508 1183 -1492 1217
rect -1458 1183 -1442 1217
rect -1508 1167 -1442 1183
rect -1390 1217 -1324 1233
rect -1390 1183 -1374 1217
rect -1340 1183 -1324 1217
rect -1390 1167 -1324 1183
rect -1272 1217 -1206 1233
rect -1272 1183 -1256 1217
rect -1222 1183 -1206 1217
rect -1272 1167 -1206 1183
rect -1154 1217 -1088 1233
rect -1154 1183 -1138 1217
rect -1104 1183 -1088 1217
rect -1154 1167 -1088 1183
rect -1036 1217 -970 1233
rect -1036 1183 -1020 1217
rect -986 1183 -970 1217
rect -1036 1167 -970 1183
rect -918 1217 -852 1233
rect -918 1183 -902 1217
rect -868 1183 -852 1217
rect -918 1167 -852 1183
rect -800 1217 -734 1233
rect -800 1183 -784 1217
rect -750 1183 -734 1217
rect -800 1167 -734 1183
rect -682 1217 -616 1233
rect -682 1183 -666 1217
rect -632 1183 -616 1217
rect -682 1167 -616 1183
rect -564 1217 -498 1233
rect -564 1183 -548 1217
rect -514 1183 -498 1217
rect -564 1167 -498 1183
rect -446 1217 -380 1233
rect -446 1183 -430 1217
rect -396 1183 -380 1217
rect -446 1167 -380 1183
rect -328 1217 -262 1233
rect -328 1183 -312 1217
rect -278 1183 -262 1217
rect -328 1167 -262 1183
rect -210 1217 -144 1233
rect -210 1183 -194 1217
rect -160 1183 -144 1217
rect -210 1167 -144 1183
rect -92 1217 -26 1233
rect -92 1183 -76 1217
rect -42 1183 -26 1217
rect -92 1167 -26 1183
rect 26 1217 92 1233
rect 26 1183 42 1217
rect 76 1183 92 1217
rect 26 1167 92 1183
rect 144 1217 210 1233
rect 144 1183 160 1217
rect 194 1183 210 1217
rect 144 1167 210 1183
rect 262 1217 328 1233
rect 262 1183 278 1217
rect 312 1183 328 1217
rect 262 1167 328 1183
rect 380 1217 446 1233
rect 380 1183 396 1217
rect 430 1183 446 1217
rect 380 1167 446 1183
rect 498 1217 564 1233
rect 498 1183 514 1217
rect 548 1183 564 1217
rect 498 1167 564 1183
rect 616 1217 682 1233
rect 616 1183 632 1217
rect 666 1183 682 1217
rect 616 1167 682 1183
rect 734 1217 800 1233
rect 734 1183 750 1217
rect 784 1183 800 1217
rect 734 1167 800 1183
rect 852 1217 918 1233
rect 852 1183 868 1217
rect 902 1183 918 1217
rect 852 1167 918 1183
rect 970 1217 1036 1233
rect 970 1183 986 1217
rect 1020 1183 1036 1217
rect 970 1167 1036 1183
rect 1088 1217 1154 1233
rect 1088 1183 1104 1217
rect 1138 1183 1154 1217
rect 1088 1167 1154 1183
rect 1206 1217 1272 1233
rect 1206 1183 1222 1217
rect 1256 1183 1272 1217
rect 1206 1167 1272 1183
rect 1324 1217 1390 1233
rect 1324 1183 1340 1217
rect 1374 1183 1390 1217
rect 1324 1167 1390 1183
rect 1442 1217 1508 1233
rect 1442 1183 1458 1217
rect 1492 1183 1508 1217
rect 1442 1167 1508 1183
rect 1560 1217 1626 1233
rect 1560 1183 1576 1217
rect 1610 1183 1626 1217
rect 1560 1167 1626 1183
rect 1678 1217 1744 1233
rect 1678 1183 1694 1217
rect 1728 1183 1744 1217
rect 1678 1167 1744 1183
rect 1796 1217 1862 1233
rect 1796 1183 1812 1217
rect 1846 1183 1862 1217
rect 1796 1167 1862 1183
rect 1914 1217 1980 1233
rect 1914 1183 1930 1217
rect 1964 1183 1980 1217
rect 1914 1167 1980 1183
rect 2032 1217 2098 1233
rect 2032 1183 2048 1217
rect 2082 1183 2098 1217
rect 2032 1167 2098 1183
rect 2150 1217 2216 1233
rect 2150 1183 2166 1217
rect 2200 1183 2216 1217
rect 2150 1167 2216 1183
rect 2268 1217 2334 1233
rect 2268 1183 2284 1217
rect 2318 1183 2334 1217
rect 2268 1167 2334 1183
rect 2386 1217 2452 1233
rect 2386 1183 2402 1217
rect 2436 1183 2452 1217
rect 2386 1167 2452 1183
rect 2504 1217 2570 1233
rect 2504 1183 2520 1217
rect 2554 1183 2570 1217
rect 2504 1167 2570 1183
rect 2622 1217 2688 1233
rect 2622 1183 2638 1217
rect 2672 1183 2688 1217
rect 2622 1167 2688 1183
rect 2740 1217 2806 1233
rect 2740 1183 2756 1217
rect 2790 1183 2806 1217
rect 2740 1167 2806 1183
rect 2858 1217 2924 1233
rect 2858 1183 2874 1217
rect 2908 1183 2924 1217
rect 2858 1167 2924 1183
rect -2921 1136 -2861 1167
rect -2803 1136 -2743 1167
rect -2685 1136 -2625 1167
rect -2567 1136 -2507 1167
rect -2449 1136 -2389 1167
rect -2331 1136 -2271 1167
rect -2213 1136 -2153 1167
rect -2095 1136 -2035 1167
rect -1977 1136 -1917 1167
rect -1859 1136 -1799 1167
rect -1741 1136 -1681 1167
rect -1623 1136 -1563 1167
rect -1505 1136 -1445 1167
rect -1387 1136 -1327 1167
rect -1269 1136 -1209 1167
rect -1151 1136 -1091 1167
rect -1033 1136 -973 1167
rect -915 1136 -855 1167
rect -797 1136 -737 1167
rect -679 1136 -619 1167
rect -561 1136 -501 1167
rect -443 1136 -383 1167
rect -325 1136 -265 1167
rect -207 1136 -147 1167
rect -89 1136 -29 1167
rect 29 1136 89 1167
rect 147 1136 207 1167
rect 265 1136 325 1167
rect 383 1136 443 1167
rect 501 1136 561 1167
rect 619 1136 679 1167
rect 737 1136 797 1167
rect 855 1136 915 1167
rect 973 1136 1033 1167
rect 1091 1136 1151 1167
rect 1209 1136 1269 1167
rect 1327 1136 1387 1167
rect 1445 1136 1505 1167
rect 1563 1136 1623 1167
rect 1681 1136 1741 1167
rect 1799 1136 1859 1167
rect 1917 1136 1977 1167
rect 2035 1136 2095 1167
rect 2153 1136 2213 1167
rect 2271 1136 2331 1167
rect 2389 1136 2449 1167
rect 2507 1136 2567 1167
rect 2625 1136 2685 1167
rect 2743 1136 2803 1167
rect 2861 1136 2921 1167
rect -2921 505 -2861 536
rect -2803 505 -2743 536
rect -2685 505 -2625 536
rect -2567 505 -2507 536
rect -2449 505 -2389 536
rect -2331 505 -2271 536
rect -2213 505 -2153 536
rect -2095 505 -2035 536
rect -1977 505 -1917 536
rect -1859 505 -1799 536
rect -1741 505 -1681 536
rect -1623 505 -1563 536
rect -1505 505 -1445 536
rect -1387 505 -1327 536
rect -1269 505 -1209 536
rect -1151 505 -1091 536
rect -1033 505 -973 536
rect -915 505 -855 536
rect -797 505 -737 536
rect -679 505 -619 536
rect -561 505 -501 536
rect -443 505 -383 536
rect -325 505 -265 536
rect -207 505 -147 536
rect -89 505 -29 536
rect 29 505 89 536
rect 147 505 207 536
rect 265 505 325 536
rect 383 505 443 536
rect 501 505 561 536
rect 619 505 679 536
rect 737 505 797 536
rect 855 505 915 536
rect 973 505 1033 536
rect 1091 505 1151 536
rect 1209 505 1269 536
rect 1327 505 1387 536
rect 1445 505 1505 536
rect 1563 505 1623 536
rect 1681 505 1741 536
rect 1799 505 1859 536
rect 1917 505 1977 536
rect 2035 505 2095 536
rect 2153 505 2213 536
rect 2271 505 2331 536
rect 2389 505 2449 536
rect 2507 505 2567 536
rect 2625 505 2685 536
rect 2743 505 2803 536
rect 2861 505 2921 536
rect -2924 489 -2858 505
rect -2924 455 -2908 489
rect -2874 455 -2858 489
rect -2924 439 -2858 455
rect -2806 489 -2740 505
rect -2806 455 -2790 489
rect -2756 455 -2740 489
rect -2806 439 -2740 455
rect -2688 489 -2622 505
rect -2688 455 -2672 489
rect -2638 455 -2622 489
rect -2688 439 -2622 455
rect -2570 489 -2504 505
rect -2570 455 -2554 489
rect -2520 455 -2504 489
rect -2570 439 -2504 455
rect -2452 489 -2386 505
rect -2452 455 -2436 489
rect -2402 455 -2386 489
rect -2452 439 -2386 455
rect -2334 489 -2268 505
rect -2334 455 -2318 489
rect -2284 455 -2268 489
rect -2334 439 -2268 455
rect -2216 489 -2150 505
rect -2216 455 -2200 489
rect -2166 455 -2150 489
rect -2216 439 -2150 455
rect -2098 489 -2032 505
rect -2098 455 -2082 489
rect -2048 455 -2032 489
rect -2098 439 -2032 455
rect -1980 489 -1914 505
rect -1980 455 -1964 489
rect -1930 455 -1914 489
rect -1980 439 -1914 455
rect -1862 489 -1796 505
rect -1862 455 -1846 489
rect -1812 455 -1796 489
rect -1862 439 -1796 455
rect -1744 489 -1678 505
rect -1744 455 -1728 489
rect -1694 455 -1678 489
rect -1744 439 -1678 455
rect -1626 489 -1560 505
rect -1626 455 -1610 489
rect -1576 455 -1560 489
rect -1626 439 -1560 455
rect -1508 489 -1442 505
rect -1508 455 -1492 489
rect -1458 455 -1442 489
rect -1508 439 -1442 455
rect -1390 489 -1324 505
rect -1390 455 -1374 489
rect -1340 455 -1324 489
rect -1390 439 -1324 455
rect -1272 489 -1206 505
rect -1272 455 -1256 489
rect -1222 455 -1206 489
rect -1272 439 -1206 455
rect -1154 489 -1088 505
rect -1154 455 -1138 489
rect -1104 455 -1088 489
rect -1154 439 -1088 455
rect -1036 489 -970 505
rect -1036 455 -1020 489
rect -986 455 -970 489
rect -1036 439 -970 455
rect -918 489 -852 505
rect -918 455 -902 489
rect -868 455 -852 489
rect -918 439 -852 455
rect -800 489 -734 505
rect -800 455 -784 489
rect -750 455 -734 489
rect -800 439 -734 455
rect -682 489 -616 505
rect -682 455 -666 489
rect -632 455 -616 489
rect -682 439 -616 455
rect -564 489 -498 505
rect -564 455 -548 489
rect -514 455 -498 489
rect -564 439 -498 455
rect -446 489 -380 505
rect -446 455 -430 489
rect -396 455 -380 489
rect -446 439 -380 455
rect -328 489 -262 505
rect -328 455 -312 489
rect -278 455 -262 489
rect -328 439 -262 455
rect -210 489 -144 505
rect -210 455 -194 489
rect -160 455 -144 489
rect -210 439 -144 455
rect -92 489 -26 505
rect -92 455 -76 489
rect -42 455 -26 489
rect -92 439 -26 455
rect 26 489 92 505
rect 26 455 42 489
rect 76 455 92 489
rect 26 439 92 455
rect 144 489 210 505
rect 144 455 160 489
rect 194 455 210 489
rect 144 439 210 455
rect 262 489 328 505
rect 262 455 278 489
rect 312 455 328 489
rect 262 439 328 455
rect 380 489 446 505
rect 380 455 396 489
rect 430 455 446 489
rect 380 439 446 455
rect 498 489 564 505
rect 498 455 514 489
rect 548 455 564 489
rect 498 439 564 455
rect 616 489 682 505
rect 616 455 632 489
rect 666 455 682 489
rect 616 439 682 455
rect 734 489 800 505
rect 734 455 750 489
rect 784 455 800 489
rect 734 439 800 455
rect 852 489 918 505
rect 852 455 868 489
rect 902 455 918 489
rect 852 439 918 455
rect 970 489 1036 505
rect 970 455 986 489
rect 1020 455 1036 489
rect 970 439 1036 455
rect 1088 489 1154 505
rect 1088 455 1104 489
rect 1138 455 1154 489
rect 1088 439 1154 455
rect 1206 489 1272 505
rect 1206 455 1222 489
rect 1256 455 1272 489
rect 1206 439 1272 455
rect 1324 489 1390 505
rect 1324 455 1340 489
rect 1374 455 1390 489
rect 1324 439 1390 455
rect 1442 489 1508 505
rect 1442 455 1458 489
rect 1492 455 1508 489
rect 1442 439 1508 455
rect 1560 489 1626 505
rect 1560 455 1576 489
rect 1610 455 1626 489
rect 1560 439 1626 455
rect 1678 489 1744 505
rect 1678 455 1694 489
rect 1728 455 1744 489
rect 1678 439 1744 455
rect 1796 489 1862 505
rect 1796 455 1812 489
rect 1846 455 1862 489
rect 1796 439 1862 455
rect 1914 489 1980 505
rect 1914 455 1930 489
rect 1964 455 1980 489
rect 1914 439 1980 455
rect 2032 489 2098 505
rect 2032 455 2048 489
rect 2082 455 2098 489
rect 2032 439 2098 455
rect 2150 489 2216 505
rect 2150 455 2166 489
rect 2200 455 2216 489
rect 2150 439 2216 455
rect 2268 489 2334 505
rect 2268 455 2284 489
rect 2318 455 2334 489
rect 2268 439 2334 455
rect 2386 489 2452 505
rect 2386 455 2402 489
rect 2436 455 2452 489
rect 2386 439 2452 455
rect 2504 489 2570 505
rect 2504 455 2520 489
rect 2554 455 2570 489
rect 2504 439 2570 455
rect 2622 489 2688 505
rect 2622 455 2638 489
rect 2672 455 2688 489
rect 2622 439 2688 455
rect 2740 489 2806 505
rect 2740 455 2756 489
rect 2790 455 2806 489
rect 2740 439 2806 455
rect 2858 489 2924 505
rect 2858 455 2874 489
rect 2908 455 2924 489
rect 2858 439 2924 455
rect -2924 381 -2858 397
rect -2924 347 -2908 381
rect -2874 347 -2858 381
rect -2924 331 -2858 347
rect -2806 381 -2740 397
rect -2806 347 -2790 381
rect -2756 347 -2740 381
rect -2806 331 -2740 347
rect -2688 381 -2622 397
rect -2688 347 -2672 381
rect -2638 347 -2622 381
rect -2688 331 -2622 347
rect -2570 381 -2504 397
rect -2570 347 -2554 381
rect -2520 347 -2504 381
rect -2570 331 -2504 347
rect -2452 381 -2386 397
rect -2452 347 -2436 381
rect -2402 347 -2386 381
rect -2452 331 -2386 347
rect -2334 381 -2268 397
rect -2334 347 -2318 381
rect -2284 347 -2268 381
rect -2334 331 -2268 347
rect -2216 381 -2150 397
rect -2216 347 -2200 381
rect -2166 347 -2150 381
rect -2216 331 -2150 347
rect -2098 381 -2032 397
rect -2098 347 -2082 381
rect -2048 347 -2032 381
rect -2098 331 -2032 347
rect -1980 381 -1914 397
rect -1980 347 -1964 381
rect -1930 347 -1914 381
rect -1980 331 -1914 347
rect -1862 381 -1796 397
rect -1862 347 -1846 381
rect -1812 347 -1796 381
rect -1862 331 -1796 347
rect -1744 381 -1678 397
rect -1744 347 -1728 381
rect -1694 347 -1678 381
rect -1744 331 -1678 347
rect -1626 381 -1560 397
rect -1626 347 -1610 381
rect -1576 347 -1560 381
rect -1626 331 -1560 347
rect -1508 381 -1442 397
rect -1508 347 -1492 381
rect -1458 347 -1442 381
rect -1508 331 -1442 347
rect -1390 381 -1324 397
rect -1390 347 -1374 381
rect -1340 347 -1324 381
rect -1390 331 -1324 347
rect -1272 381 -1206 397
rect -1272 347 -1256 381
rect -1222 347 -1206 381
rect -1272 331 -1206 347
rect -1154 381 -1088 397
rect -1154 347 -1138 381
rect -1104 347 -1088 381
rect -1154 331 -1088 347
rect -1036 381 -970 397
rect -1036 347 -1020 381
rect -986 347 -970 381
rect -1036 331 -970 347
rect -918 381 -852 397
rect -918 347 -902 381
rect -868 347 -852 381
rect -918 331 -852 347
rect -800 381 -734 397
rect -800 347 -784 381
rect -750 347 -734 381
rect -800 331 -734 347
rect -682 381 -616 397
rect -682 347 -666 381
rect -632 347 -616 381
rect -682 331 -616 347
rect -564 381 -498 397
rect -564 347 -548 381
rect -514 347 -498 381
rect -564 331 -498 347
rect -446 381 -380 397
rect -446 347 -430 381
rect -396 347 -380 381
rect -446 331 -380 347
rect -328 381 -262 397
rect -328 347 -312 381
rect -278 347 -262 381
rect -328 331 -262 347
rect -210 381 -144 397
rect -210 347 -194 381
rect -160 347 -144 381
rect -210 331 -144 347
rect -92 381 -26 397
rect -92 347 -76 381
rect -42 347 -26 381
rect -92 331 -26 347
rect 26 381 92 397
rect 26 347 42 381
rect 76 347 92 381
rect 26 331 92 347
rect 144 381 210 397
rect 144 347 160 381
rect 194 347 210 381
rect 144 331 210 347
rect 262 381 328 397
rect 262 347 278 381
rect 312 347 328 381
rect 262 331 328 347
rect 380 381 446 397
rect 380 347 396 381
rect 430 347 446 381
rect 380 331 446 347
rect 498 381 564 397
rect 498 347 514 381
rect 548 347 564 381
rect 498 331 564 347
rect 616 381 682 397
rect 616 347 632 381
rect 666 347 682 381
rect 616 331 682 347
rect 734 381 800 397
rect 734 347 750 381
rect 784 347 800 381
rect 734 331 800 347
rect 852 381 918 397
rect 852 347 868 381
rect 902 347 918 381
rect 852 331 918 347
rect 970 381 1036 397
rect 970 347 986 381
rect 1020 347 1036 381
rect 970 331 1036 347
rect 1088 381 1154 397
rect 1088 347 1104 381
rect 1138 347 1154 381
rect 1088 331 1154 347
rect 1206 381 1272 397
rect 1206 347 1222 381
rect 1256 347 1272 381
rect 1206 331 1272 347
rect 1324 381 1390 397
rect 1324 347 1340 381
rect 1374 347 1390 381
rect 1324 331 1390 347
rect 1442 381 1508 397
rect 1442 347 1458 381
rect 1492 347 1508 381
rect 1442 331 1508 347
rect 1560 381 1626 397
rect 1560 347 1576 381
rect 1610 347 1626 381
rect 1560 331 1626 347
rect 1678 381 1744 397
rect 1678 347 1694 381
rect 1728 347 1744 381
rect 1678 331 1744 347
rect 1796 381 1862 397
rect 1796 347 1812 381
rect 1846 347 1862 381
rect 1796 331 1862 347
rect 1914 381 1980 397
rect 1914 347 1930 381
rect 1964 347 1980 381
rect 1914 331 1980 347
rect 2032 381 2098 397
rect 2032 347 2048 381
rect 2082 347 2098 381
rect 2032 331 2098 347
rect 2150 381 2216 397
rect 2150 347 2166 381
rect 2200 347 2216 381
rect 2150 331 2216 347
rect 2268 381 2334 397
rect 2268 347 2284 381
rect 2318 347 2334 381
rect 2268 331 2334 347
rect 2386 381 2452 397
rect 2386 347 2402 381
rect 2436 347 2452 381
rect 2386 331 2452 347
rect 2504 381 2570 397
rect 2504 347 2520 381
rect 2554 347 2570 381
rect 2504 331 2570 347
rect 2622 381 2688 397
rect 2622 347 2638 381
rect 2672 347 2688 381
rect 2622 331 2688 347
rect 2740 381 2806 397
rect 2740 347 2756 381
rect 2790 347 2806 381
rect 2740 331 2806 347
rect 2858 381 2924 397
rect 2858 347 2874 381
rect 2908 347 2924 381
rect 2858 331 2924 347
rect -2921 300 -2861 331
rect -2803 300 -2743 331
rect -2685 300 -2625 331
rect -2567 300 -2507 331
rect -2449 300 -2389 331
rect -2331 300 -2271 331
rect -2213 300 -2153 331
rect -2095 300 -2035 331
rect -1977 300 -1917 331
rect -1859 300 -1799 331
rect -1741 300 -1681 331
rect -1623 300 -1563 331
rect -1505 300 -1445 331
rect -1387 300 -1327 331
rect -1269 300 -1209 331
rect -1151 300 -1091 331
rect -1033 300 -973 331
rect -915 300 -855 331
rect -797 300 -737 331
rect -679 300 -619 331
rect -561 300 -501 331
rect -443 300 -383 331
rect -325 300 -265 331
rect -207 300 -147 331
rect -89 300 -29 331
rect 29 300 89 331
rect 147 300 207 331
rect 265 300 325 331
rect 383 300 443 331
rect 501 300 561 331
rect 619 300 679 331
rect 737 300 797 331
rect 855 300 915 331
rect 973 300 1033 331
rect 1091 300 1151 331
rect 1209 300 1269 331
rect 1327 300 1387 331
rect 1445 300 1505 331
rect 1563 300 1623 331
rect 1681 300 1741 331
rect 1799 300 1859 331
rect 1917 300 1977 331
rect 2035 300 2095 331
rect 2153 300 2213 331
rect 2271 300 2331 331
rect 2389 300 2449 331
rect 2507 300 2567 331
rect 2625 300 2685 331
rect 2743 300 2803 331
rect 2861 300 2921 331
rect -2921 -331 -2861 -300
rect -2803 -331 -2743 -300
rect -2685 -331 -2625 -300
rect -2567 -331 -2507 -300
rect -2449 -331 -2389 -300
rect -2331 -331 -2271 -300
rect -2213 -331 -2153 -300
rect -2095 -331 -2035 -300
rect -1977 -331 -1917 -300
rect -1859 -331 -1799 -300
rect -1741 -331 -1681 -300
rect -1623 -331 -1563 -300
rect -1505 -331 -1445 -300
rect -1387 -331 -1327 -300
rect -1269 -331 -1209 -300
rect -1151 -331 -1091 -300
rect -1033 -331 -973 -300
rect -915 -331 -855 -300
rect -797 -331 -737 -300
rect -679 -331 -619 -300
rect -561 -331 -501 -300
rect -443 -331 -383 -300
rect -325 -331 -265 -300
rect -207 -331 -147 -300
rect -89 -331 -29 -300
rect 29 -331 89 -300
rect 147 -331 207 -300
rect 265 -331 325 -300
rect 383 -331 443 -300
rect 501 -331 561 -300
rect 619 -331 679 -300
rect 737 -331 797 -300
rect 855 -331 915 -300
rect 973 -331 1033 -300
rect 1091 -331 1151 -300
rect 1209 -331 1269 -300
rect 1327 -331 1387 -300
rect 1445 -331 1505 -300
rect 1563 -331 1623 -300
rect 1681 -331 1741 -300
rect 1799 -331 1859 -300
rect 1917 -331 1977 -300
rect 2035 -331 2095 -300
rect 2153 -331 2213 -300
rect 2271 -331 2331 -300
rect 2389 -331 2449 -300
rect 2507 -331 2567 -300
rect 2625 -331 2685 -300
rect 2743 -331 2803 -300
rect 2861 -331 2921 -300
rect -2924 -347 -2858 -331
rect -2924 -381 -2908 -347
rect -2874 -381 -2858 -347
rect -2924 -397 -2858 -381
rect -2806 -347 -2740 -331
rect -2806 -381 -2790 -347
rect -2756 -381 -2740 -347
rect -2806 -397 -2740 -381
rect -2688 -347 -2622 -331
rect -2688 -381 -2672 -347
rect -2638 -381 -2622 -347
rect -2688 -397 -2622 -381
rect -2570 -347 -2504 -331
rect -2570 -381 -2554 -347
rect -2520 -381 -2504 -347
rect -2570 -397 -2504 -381
rect -2452 -347 -2386 -331
rect -2452 -381 -2436 -347
rect -2402 -381 -2386 -347
rect -2452 -397 -2386 -381
rect -2334 -347 -2268 -331
rect -2334 -381 -2318 -347
rect -2284 -381 -2268 -347
rect -2334 -397 -2268 -381
rect -2216 -347 -2150 -331
rect -2216 -381 -2200 -347
rect -2166 -381 -2150 -347
rect -2216 -397 -2150 -381
rect -2098 -347 -2032 -331
rect -2098 -381 -2082 -347
rect -2048 -381 -2032 -347
rect -2098 -397 -2032 -381
rect -1980 -347 -1914 -331
rect -1980 -381 -1964 -347
rect -1930 -381 -1914 -347
rect -1980 -397 -1914 -381
rect -1862 -347 -1796 -331
rect -1862 -381 -1846 -347
rect -1812 -381 -1796 -347
rect -1862 -397 -1796 -381
rect -1744 -347 -1678 -331
rect -1744 -381 -1728 -347
rect -1694 -381 -1678 -347
rect -1744 -397 -1678 -381
rect -1626 -347 -1560 -331
rect -1626 -381 -1610 -347
rect -1576 -381 -1560 -347
rect -1626 -397 -1560 -381
rect -1508 -347 -1442 -331
rect -1508 -381 -1492 -347
rect -1458 -381 -1442 -347
rect -1508 -397 -1442 -381
rect -1390 -347 -1324 -331
rect -1390 -381 -1374 -347
rect -1340 -381 -1324 -347
rect -1390 -397 -1324 -381
rect -1272 -347 -1206 -331
rect -1272 -381 -1256 -347
rect -1222 -381 -1206 -347
rect -1272 -397 -1206 -381
rect -1154 -347 -1088 -331
rect -1154 -381 -1138 -347
rect -1104 -381 -1088 -347
rect -1154 -397 -1088 -381
rect -1036 -347 -970 -331
rect -1036 -381 -1020 -347
rect -986 -381 -970 -347
rect -1036 -397 -970 -381
rect -918 -347 -852 -331
rect -918 -381 -902 -347
rect -868 -381 -852 -347
rect -918 -397 -852 -381
rect -800 -347 -734 -331
rect -800 -381 -784 -347
rect -750 -381 -734 -347
rect -800 -397 -734 -381
rect -682 -347 -616 -331
rect -682 -381 -666 -347
rect -632 -381 -616 -347
rect -682 -397 -616 -381
rect -564 -347 -498 -331
rect -564 -381 -548 -347
rect -514 -381 -498 -347
rect -564 -397 -498 -381
rect -446 -347 -380 -331
rect -446 -381 -430 -347
rect -396 -381 -380 -347
rect -446 -397 -380 -381
rect -328 -347 -262 -331
rect -328 -381 -312 -347
rect -278 -381 -262 -347
rect -328 -397 -262 -381
rect -210 -347 -144 -331
rect -210 -381 -194 -347
rect -160 -381 -144 -347
rect -210 -397 -144 -381
rect -92 -347 -26 -331
rect -92 -381 -76 -347
rect -42 -381 -26 -347
rect -92 -397 -26 -381
rect 26 -347 92 -331
rect 26 -381 42 -347
rect 76 -381 92 -347
rect 26 -397 92 -381
rect 144 -347 210 -331
rect 144 -381 160 -347
rect 194 -381 210 -347
rect 144 -397 210 -381
rect 262 -347 328 -331
rect 262 -381 278 -347
rect 312 -381 328 -347
rect 262 -397 328 -381
rect 380 -347 446 -331
rect 380 -381 396 -347
rect 430 -381 446 -347
rect 380 -397 446 -381
rect 498 -347 564 -331
rect 498 -381 514 -347
rect 548 -381 564 -347
rect 498 -397 564 -381
rect 616 -347 682 -331
rect 616 -381 632 -347
rect 666 -381 682 -347
rect 616 -397 682 -381
rect 734 -347 800 -331
rect 734 -381 750 -347
rect 784 -381 800 -347
rect 734 -397 800 -381
rect 852 -347 918 -331
rect 852 -381 868 -347
rect 902 -381 918 -347
rect 852 -397 918 -381
rect 970 -347 1036 -331
rect 970 -381 986 -347
rect 1020 -381 1036 -347
rect 970 -397 1036 -381
rect 1088 -347 1154 -331
rect 1088 -381 1104 -347
rect 1138 -381 1154 -347
rect 1088 -397 1154 -381
rect 1206 -347 1272 -331
rect 1206 -381 1222 -347
rect 1256 -381 1272 -347
rect 1206 -397 1272 -381
rect 1324 -347 1390 -331
rect 1324 -381 1340 -347
rect 1374 -381 1390 -347
rect 1324 -397 1390 -381
rect 1442 -347 1508 -331
rect 1442 -381 1458 -347
rect 1492 -381 1508 -347
rect 1442 -397 1508 -381
rect 1560 -347 1626 -331
rect 1560 -381 1576 -347
rect 1610 -381 1626 -347
rect 1560 -397 1626 -381
rect 1678 -347 1744 -331
rect 1678 -381 1694 -347
rect 1728 -381 1744 -347
rect 1678 -397 1744 -381
rect 1796 -347 1862 -331
rect 1796 -381 1812 -347
rect 1846 -381 1862 -347
rect 1796 -397 1862 -381
rect 1914 -347 1980 -331
rect 1914 -381 1930 -347
rect 1964 -381 1980 -347
rect 1914 -397 1980 -381
rect 2032 -347 2098 -331
rect 2032 -381 2048 -347
rect 2082 -381 2098 -347
rect 2032 -397 2098 -381
rect 2150 -347 2216 -331
rect 2150 -381 2166 -347
rect 2200 -381 2216 -347
rect 2150 -397 2216 -381
rect 2268 -347 2334 -331
rect 2268 -381 2284 -347
rect 2318 -381 2334 -347
rect 2268 -397 2334 -381
rect 2386 -347 2452 -331
rect 2386 -381 2402 -347
rect 2436 -381 2452 -347
rect 2386 -397 2452 -381
rect 2504 -347 2570 -331
rect 2504 -381 2520 -347
rect 2554 -381 2570 -347
rect 2504 -397 2570 -381
rect 2622 -347 2688 -331
rect 2622 -381 2638 -347
rect 2672 -381 2688 -347
rect 2622 -397 2688 -381
rect 2740 -347 2806 -331
rect 2740 -381 2756 -347
rect 2790 -381 2806 -347
rect 2740 -397 2806 -381
rect 2858 -347 2924 -331
rect 2858 -381 2874 -347
rect 2908 -381 2924 -347
rect 2858 -397 2924 -381
rect -2924 -455 -2858 -439
rect -2924 -489 -2908 -455
rect -2874 -489 -2858 -455
rect -2924 -505 -2858 -489
rect -2806 -455 -2740 -439
rect -2806 -489 -2790 -455
rect -2756 -489 -2740 -455
rect -2806 -505 -2740 -489
rect -2688 -455 -2622 -439
rect -2688 -489 -2672 -455
rect -2638 -489 -2622 -455
rect -2688 -505 -2622 -489
rect -2570 -455 -2504 -439
rect -2570 -489 -2554 -455
rect -2520 -489 -2504 -455
rect -2570 -505 -2504 -489
rect -2452 -455 -2386 -439
rect -2452 -489 -2436 -455
rect -2402 -489 -2386 -455
rect -2452 -505 -2386 -489
rect -2334 -455 -2268 -439
rect -2334 -489 -2318 -455
rect -2284 -489 -2268 -455
rect -2334 -505 -2268 -489
rect -2216 -455 -2150 -439
rect -2216 -489 -2200 -455
rect -2166 -489 -2150 -455
rect -2216 -505 -2150 -489
rect -2098 -455 -2032 -439
rect -2098 -489 -2082 -455
rect -2048 -489 -2032 -455
rect -2098 -505 -2032 -489
rect -1980 -455 -1914 -439
rect -1980 -489 -1964 -455
rect -1930 -489 -1914 -455
rect -1980 -505 -1914 -489
rect -1862 -455 -1796 -439
rect -1862 -489 -1846 -455
rect -1812 -489 -1796 -455
rect -1862 -505 -1796 -489
rect -1744 -455 -1678 -439
rect -1744 -489 -1728 -455
rect -1694 -489 -1678 -455
rect -1744 -505 -1678 -489
rect -1626 -455 -1560 -439
rect -1626 -489 -1610 -455
rect -1576 -489 -1560 -455
rect -1626 -505 -1560 -489
rect -1508 -455 -1442 -439
rect -1508 -489 -1492 -455
rect -1458 -489 -1442 -455
rect -1508 -505 -1442 -489
rect -1390 -455 -1324 -439
rect -1390 -489 -1374 -455
rect -1340 -489 -1324 -455
rect -1390 -505 -1324 -489
rect -1272 -455 -1206 -439
rect -1272 -489 -1256 -455
rect -1222 -489 -1206 -455
rect -1272 -505 -1206 -489
rect -1154 -455 -1088 -439
rect -1154 -489 -1138 -455
rect -1104 -489 -1088 -455
rect -1154 -505 -1088 -489
rect -1036 -455 -970 -439
rect -1036 -489 -1020 -455
rect -986 -489 -970 -455
rect -1036 -505 -970 -489
rect -918 -455 -852 -439
rect -918 -489 -902 -455
rect -868 -489 -852 -455
rect -918 -505 -852 -489
rect -800 -455 -734 -439
rect -800 -489 -784 -455
rect -750 -489 -734 -455
rect -800 -505 -734 -489
rect -682 -455 -616 -439
rect -682 -489 -666 -455
rect -632 -489 -616 -455
rect -682 -505 -616 -489
rect -564 -455 -498 -439
rect -564 -489 -548 -455
rect -514 -489 -498 -455
rect -564 -505 -498 -489
rect -446 -455 -380 -439
rect -446 -489 -430 -455
rect -396 -489 -380 -455
rect -446 -505 -380 -489
rect -328 -455 -262 -439
rect -328 -489 -312 -455
rect -278 -489 -262 -455
rect -328 -505 -262 -489
rect -210 -455 -144 -439
rect -210 -489 -194 -455
rect -160 -489 -144 -455
rect -210 -505 -144 -489
rect -92 -455 -26 -439
rect -92 -489 -76 -455
rect -42 -489 -26 -455
rect -92 -505 -26 -489
rect 26 -455 92 -439
rect 26 -489 42 -455
rect 76 -489 92 -455
rect 26 -505 92 -489
rect 144 -455 210 -439
rect 144 -489 160 -455
rect 194 -489 210 -455
rect 144 -505 210 -489
rect 262 -455 328 -439
rect 262 -489 278 -455
rect 312 -489 328 -455
rect 262 -505 328 -489
rect 380 -455 446 -439
rect 380 -489 396 -455
rect 430 -489 446 -455
rect 380 -505 446 -489
rect 498 -455 564 -439
rect 498 -489 514 -455
rect 548 -489 564 -455
rect 498 -505 564 -489
rect 616 -455 682 -439
rect 616 -489 632 -455
rect 666 -489 682 -455
rect 616 -505 682 -489
rect 734 -455 800 -439
rect 734 -489 750 -455
rect 784 -489 800 -455
rect 734 -505 800 -489
rect 852 -455 918 -439
rect 852 -489 868 -455
rect 902 -489 918 -455
rect 852 -505 918 -489
rect 970 -455 1036 -439
rect 970 -489 986 -455
rect 1020 -489 1036 -455
rect 970 -505 1036 -489
rect 1088 -455 1154 -439
rect 1088 -489 1104 -455
rect 1138 -489 1154 -455
rect 1088 -505 1154 -489
rect 1206 -455 1272 -439
rect 1206 -489 1222 -455
rect 1256 -489 1272 -455
rect 1206 -505 1272 -489
rect 1324 -455 1390 -439
rect 1324 -489 1340 -455
rect 1374 -489 1390 -455
rect 1324 -505 1390 -489
rect 1442 -455 1508 -439
rect 1442 -489 1458 -455
rect 1492 -489 1508 -455
rect 1442 -505 1508 -489
rect 1560 -455 1626 -439
rect 1560 -489 1576 -455
rect 1610 -489 1626 -455
rect 1560 -505 1626 -489
rect 1678 -455 1744 -439
rect 1678 -489 1694 -455
rect 1728 -489 1744 -455
rect 1678 -505 1744 -489
rect 1796 -455 1862 -439
rect 1796 -489 1812 -455
rect 1846 -489 1862 -455
rect 1796 -505 1862 -489
rect 1914 -455 1980 -439
rect 1914 -489 1930 -455
rect 1964 -489 1980 -455
rect 1914 -505 1980 -489
rect 2032 -455 2098 -439
rect 2032 -489 2048 -455
rect 2082 -489 2098 -455
rect 2032 -505 2098 -489
rect 2150 -455 2216 -439
rect 2150 -489 2166 -455
rect 2200 -489 2216 -455
rect 2150 -505 2216 -489
rect 2268 -455 2334 -439
rect 2268 -489 2284 -455
rect 2318 -489 2334 -455
rect 2268 -505 2334 -489
rect 2386 -455 2452 -439
rect 2386 -489 2402 -455
rect 2436 -489 2452 -455
rect 2386 -505 2452 -489
rect 2504 -455 2570 -439
rect 2504 -489 2520 -455
rect 2554 -489 2570 -455
rect 2504 -505 2570 -489
rect 2622 -455 2688 -439
rect 2622 -489 2638 -455
rect 2672 -489 2688 -455
rect 2622 -505 2688 -489
rect 2740 -455 2806 -439
rect 2740 -489 2756 -455
rect 2790 -489 2806 -455
rect 2740 -505 2806 -489
rect 2858 -455 2924 -439
rect 2858 -489 2874 -455
rect 2908 -489 2924 -455
rect 2858 -505 2924 -489
rect -2921 -536 -2861 -505
rect -2803 -536 -2743 -505
rect -2685 -536 -2625 -505
rect -2567 -536 -2507 -505
rect -2449 -536 -2389 -505
rect -2331 -536 -2271 -505
rect -2213 -536 -2153 -505
rect -2095 -536 -2035 -505
rect -1977 -536 -1917 -505
rect -1859 -536 -1799 -505
rect -1741 -536 -1681 -505
rect -1623 -536 -1563 -505
rect -1505 -536 -1445 -505
rect -1387 -536 -1327 -505
rect -1269 -536 -1209 -505
rect -1151 -536 -1091 -505
rect -1033 -536 -973 -505
rect -915 -536 -855 -505
rect -797 -536 -737 -505
rect -679 -536 -619 -505
rect -561 -536 -501 -505
rect -443 -536 -383 -505
rect -325 -536 -265 -505
rect -207 -536 -147 -505
rect -89 -536 -29 -505
rect 29 -536 89 -505
rect 147 -536 207 -505
rect 265 -536 325 -505
rect 383 -536 443 -505
rect 501 -536 561 -505
rect 619 -536 679 -505
rect 737 -536 797 -505
rect 855 -536 915 -505
rect 973 -536 1033 -505
rect 1091 -536 1151 -505
rect 1209 -536 1269 -505
rect 1327 -536 1387 -505
rect 1445 -536 1505 -505
rect 1563 -536 1623 -505
rect 1681 -536 1741 -505
rect 1799 -536 1859 -505
rect 1917 -536 1977 -505
rect 2035 -536 2095 -505
rect 2153 -536 2213 -505
rect 2271 -536 2331 -505
rect 2389 -536 2449 -505
rect 2507 -536 2567 -505
rect 2625 -536 2685 -505
rect 2743 -536 2803 -505
rect 2861 -536 2921 -505
rect -2921 -1167 -2861 -1136
rect -2803 -1167 -2743 -1136
rect -2685 -1167 -2625 -1136
rect -2567 -1167 -2507 -1136
rect -2449 -1167 -2389 -1136
rect -2331 -1167 -2271 -1136
rect -2213 -1167 -2153 -1136
rect -2095 -1167 -2035 -1136
rect -1977 -1167 -1917 -1136
rect -1859 -1167 -1799 -1136
rect -1741 -1167 -1681 -1136
rect -1623 -1167 -1563 -1136
rect -1505 -1167 -1445 -1136
rect -1387 -1167 -1327 -1136
rect -1269 -1167 -1209 -1136
rect -1151 -1167 -1091 -1136
rect -1033 -1167 -973 -1136
rect -915 -1167 -855 -1136
rect -797 -1167 -737 -1136
rect -679 -1167 -619 -1136
rect -561 -1167 -501 -1136
rect -443 -1167 -383 -1136
rect -325 -1167 -265 -1136
rect -207 -1167 -147 -1136
rect -89 -1167 -29 -1136
rect 29 -1167 89 -1136
rect 147 -1167 207 -1136
rect 265 -1167 325 -1136
rect 383 -1167 443 -1136
rect 501 -1167 561 -1136
rect 619 -1167 679 -1136
rect 737 -1167 797 -1136
rect 855 -1167 915 -1136
rect 973 -1167 1033 -1136
rect 1091 -1167 1151 -1136
rect 1209 -1167 1269 -1136
rect 1327 -1167 1387 -1136
rect 1445 -1167 1505 -1136
rect 1563 -1167 1623 -1136
rect 1681 -1167 1741 -1136
rect 1799 -1167 1859 -1136
rect 1917 -1167 1977 -1136
rect 2035 -1167 2095 -1136
rect 2153 -1167 2213 -1136
rect 2271 -1167 2331 -1136
rect 2389 -1167 2449 -1136
rect 2507 -1167 2567 -1136
rect 2625 -1167 2685 -1136
rect 2743 -1167 2803 -1136
rect 2861 -1167 2921 -1136
rect -2924 -1183 -2858 -1167
rect -2924 -1217 -2908 -1183
rect -2874 -1217 -2858 -1183
rect -2924 -1233 -2858 -1217
rect -2806 -1183 -2740 -1167
rect -2806 -1217 -2790 -1183
rect -2756 -1217 -2740 -1183
rect -2806 -1233 -2740 -1217
rect -2688 -1183 -2622 -1167
rect -2688 -1217 -2672 -1183
rect -2638 -1217 -2622 -1183
rect -2688 -1233 -2622 -1217
rect -2570 -1183 -2504 -1167
rect -2570 -1217 -2554 -1183
rect -2520 -1217 -2504 -1183
rect -2570 -1233 -2504 -1217
rect -2452 -1183 -2386 -1167
rect -2452 -1217 -2436 -1183
rect -2402 -1217 -2386 -1183
rect -2452 -1233 -2386 -1217
rect -2334 -1183 -2268 -1167
rect -2334 -1217 -2318 -1183
rect -2284 -1217 -2268 -1183
rect -2334 -1233 -2268 -1217
rect -2216 -1183 -2150 -1167
rect -2216 -1217 -2200 -1183
rect -2166 -1217 -2150 -1183
rect -2216 -1233 -2150 -1217
rect -2098 -1183 -2032 -1167
rect -2098 -1217 -2082 -1183
rect -2048 -1217 -2032 -1183
rect -2098 -1233 -2032 -1217
rect -1980 -1183 -1914 -1167
rect -1980 -1217 -1964 -1183
rect -1930 -1217 -1914 -1183
rect -1980 -1233 -1914 -1217
rect -1862 -1183 -1796 -1167
rect -1862 -1217 -1846 -1183
rect -1812 -1217 -1796 -1183
rect -1862 -1233 -1796 -1217
rect -1744 -1183 -1678 -1167
rect -1744 -1217 -1728 -1183
rect -1694 -1217 -1678 -1183
rect -1744 -1233 -1678 -1217
rect -1626 -1183 -1560 -1167
rect -1626 -1217 -1610 -1183
rect -1576 -1217 -1560 -1183
rect -1626 -1233 -1560 -1217
rect -1508 -1183 -1442 -1167
rect -1508 -1217 -1492 -1183
rect -1458 -1217 -1442 -1183
rect -1508 -1233 -1442 -1217
rect -1390 -1183 -1324 -1167
rect -1390 -1217 -1374 -1183
rect -1340 -1217 -1324 -1183
rect -1390 -1233 -1324 -1217
rect -1272 -1183 -1206 -1167
rect -1272 -1217 -1256 -1183
rect -1222 -1217 -1206 -1183
rect -1272 -1233 -1206 -1217
rect -1154 -1183 -1088 -1167
rect -1154 -1217 -1138 -1183
rect -1104 -1217 -1088 -1183
rect -1154 -1233 -1088 -1217
rect -1036 -1183 -970 -1167
rect -1036 -1217 -1020 -1183
rect -986 -1217 -970 -1183
rect -1036 -1233 -970 -1217
rect -918 -1183 -852 -1167
rect -918 -1217 -902 -1183
rect -868 -1217 -852 -1183
rect -918 -1233 -852 -1217
rect -800 -1183 -734 -1167
rect -800 -1217 -784 -1183
rect -750 -1217 -734 -1183
rect -800 -1233 -734 -1217
rect -682 -1183 -616 -1167
rect -682 -1217 -666 -1183
rect -632 -1217 -616 -1183
rect -682 -1233 -616 -1217
rect -564 -1183 -498 -1167
rect -564 -1217 -548 -1183
rect -514 -1217 -498 -1183
rect -564 -1233 -498 -1217
rect -446 -1183 -380 -1167
rect -446 -1217 -430 -1183
rect -396 -1217 -380 -1183
rect -446 -1233 -380 -1217
rect -328 -1183 -262 -1167
rect -328 -1217 -312 -1183
rect -278 -1217 -262 -1183
rect -328 -1233 -262 -1217
rect -210 -1183 -144 -1167
rect -210 -1217 -194 -1183
rect -160 -1217 -144 -1183
rect -210 -1233 -144 -1217
rect -92 -1183 -26 -1167
rect -92 -1217 -76 -1183
rect -42 -1217 -26 -1183
rect -92 -1233 -26 -1217
rect 26 -1183 92 -1167
rect 26 -1217 42 -1183
rect 76 -1217 92 -1183
rect 26 -1233 92 -1217
rect 144 -1183 210 -1167
rect 144 -1217 160 -1183
rect 194 -1217 210 -1183
rect 144 -1233 210 -1217
rect 262 -1183 328 -1167
rect 262 -1217 278 -1183
rect 312 -1217 328 -1183
rect 262 -1233 328 -1217
rect 380 -1183 446 -1167
rect 380 -1217 396 -1183
rect 430 -1217 446 -1183
rect 380 -1233 446 -1217
rect 498 -1183 564 -1167
rect 498 -1217 514 -1183
rect 548 -1217 564 -1183
rect 498 -1233 564 -1217
rect 616 -1183 682 -1167
rect 616 -1217 632 -1183
rect 666 -1217 682 -1183
rect 616 -1233 682 -1217
rect 734 -1183 800 -1167
rect 734 -1217 750 -1183
rect 784 -1217 800 -1183
rect 734 -1233 800 -1217
rect 852 -1183 918 -1167
rect 852 -1217 868 -1183
rect 902 -1217 918 -1183
rect 852 -1233 918 -1217
rect 970 -1183 1036 -1167
rect 970 -1217 986 -1183
rect 1020 -1217 1036 -1183
rect 970 -1233 1036 -1217
rect 1088 -1183 1154 -1167
rect 1088 -1217 1104 -1183
rect 1138 -1217 1154 -1183
rect 1088 -1233 1154 -1217
rect 1206 -1183 1272 -1167
rect 1206 -1217 1222 -1183
rect 1256 -1217 1272 -1183
rect 1206 -1233 1272 -1217
rect 1324 -1183 1390 -1167
rect 1324 -1217 1340 -1183
rect 1374 -1217 1390 -1183
rect 1324 -1233 1390 -1217
rect 1442 -1183 1508 -1167
rect 1442 -1217 1458 -1183
rect 1492 -1217 1508 -1183
rect 1442 -1233 1508 -1217
rect 1560 -1183 1626 -1167
rect 1560 -1217 1576 -1183
rect 1610 -1217 1626 -1183
rect 1560 -1233 1626 -1217
rect 1678 -1183 1744 -1167
rect 1678 -1217 1694 -1183
rect 1728 -1217 1744 -1183
rect 1678 -1233 1744 -1217
rect 1796 -1183 1862 -1167
rect 1796 -1217 1812 -1183
rect 1846 -1217 1862 -1183
rect 1796 -1233 1862 -1217
rect 1914 -1183 1980 -1167
rect 1914 -1217 1930 -1183
rect 1964 -1217 1980 -1183
rect 1914 -1233 1980 -1217
rect 2032 -1183 2098 -1167
rect 2032 -1217 2048 -1183
rect 2082 -1217 2098 -1183
rect 2032 -1233 2098 -1217
rect 2150 -1183 2216 -1167
rect 2150 -1217 2166 -1183
rect 2200 -1217 2216 -1183
rect 2150 -1233 2216 -1217
rect 2268 -1183 2334 -1167
rect 2268 -1217 2284 -1183
rect 2318 -1217 2334 -1183
rect 2268 -1233 2334 -1217
rect 2386 -1183 2452 -1167
rect 2386 -1217 2402 -1183
rect 2436 -1217 2452 -1183
rect 2386 -1233 2452 -1217
rect 2504 -1183 2570 -1167
rect 2504 -1217 2520 -1183
rect 2554 -1217 2570 -1183
rect 2504 -1233 2570 -1217
rect 2622 -1183 2688 -1167
rect 2622 -1217 2638 -1183
rect 2672 -1217 2688 -1183
rect 2622 -1233 2688 -1217
rect 2740 -1183 2806 -1167
rect 2740 -1217 2756 -1183
rect 2790 -1217 2806 -1183
rect 2740 -1233 2806 -1217
rect 2858 -1183 2924 -1167
rect 2858 -1217 2874 -1183
rect 2908 -1217 2924 -1183
rect 2858 -1233 2924 -1217
<< polycont >>
rect -2908 1183 -2874 1217
rect -2790 1183 -2756 1217
rect -2672 1183 -2638 1217
rect -2554 1183 -2520 1217
rect -2436 1183 -2402 1217
rect -2318 1183 -2284 1217
rect -2200 1183 -2166 1217
rect -2082 1183 -2048 1217
rect -1964 1183 -1930 1217
rect -1846 1183 -1812 1217
rect -1728 1183 -1694 1217
rect -1610 1183 -1576 1217
rect -1492 1183 -1458 1217
rect -1374 1183 -1340 1217
rect -1256 1183 -1222 1217
rect -1138 1183 -1104 1217
rect -1020 1183 -986 1217
rect -902 1183 -868 1217
rect -784 1183 -750 1217
rect -666 1183 -632 1217
rect -548 1183 -514 1217
rect -430 1183 -396 1217
rect -312 1183 -278 1217
rect -194 1183 -160 1217
rect -76 1183 -42 1217
rect 42 1183 76 1217
rect 160 1183 194 1217
rect 278 1183 312 1217
rect 396 1183 430 1217
rect 514 1183 548 1217
rect 632 1183 666 1217
rect 750 1183 784 1217
rect 868 1183 902 1217
rect 986 1183 1020 1217
rect 1104 1183 1138 1217
rect 1222 1183 1256 1217
rect 1340 1183 1374 1217
rect 1458 1183 1492 1217
rect 1576 1183 1610 1217
rect 1694 1183 1728 1217
rect 1812 1183 1846 1217
rect 1930 1183 1964 1217
rect 2048 1183 2082 1217
rect 2166 1183 2200 1217
rect 2284 1183 2318 1217
rect 2402 1183 2436 1217
rect 2520 1183 2554 1217
rect 2638 1183 2672 1217
rect 2756 1183 2790 1217
rect 2874 1183 2908 1217
rect -2908 455 -2874 489
rect -2790 455 -2756 489
rect -2672 455 -2638 489
rect -2554 455 -2520 489
rect -2436 455 -2402 489
rect -2318 455 -2284 489
rect -2200 455 -2166 489
rect -2082 455 -2048 489
rect -1964 455 -1930 489
rect -1846 455 -1812 489
rect -1728 455 -1694 489
rect -1610 455 -1576 489
rect -1492 455 -1458 489
rect -1374 455 -1340 489
rect -1256 455 -1222 489
rect -1138 455 -1104 489
rect -1020 455 -986 489
rect -902 455 -868 489
rect -784 455 -750 489
rect -666 455 -632 489
rect -548 455 -514 489
rect -430 455 -396 489
rect -312 455 -278 489
rect -194 455 -160 489
rect -76 455 -42 489
rect 42 455 76 489
rect 160 455 194 489
rect 278 455 312 489
rect 396 455 430 489
rect 514 455 548 489
rect 632 455 666 489
rect 750 455 784 489
rect 868 455 902 489
rect 986 455 1020 489
rect 1104 455 1138 489
rect 1222 455 1256 489
rect 1340 455 1374 489
rect 1458 455 1492 489
rect 1576 455 1610 489
rect 1694 455 1728 489
rect 1812 455 1846 489
rect 1930 455 1964 489
rect 2048 455 2082 489
rect 2166 455 2200 489
rect 2284 455 2318 489
rect 2402 455 2436 489
rect 2520 455 2554 489
rect 2638 455 2672 489
rect 2756 455 2790 489
rect 2874 455 2908 489
rect -2908 347 -2874 381
rect -2790 347 -2756 381
rect -2672 347 -2638 381
rect -2554 347 -2520 381
rect -2436 347 -2402 381
rect -2318 347 -2284 381
rect -2200 347 -2166 381
rect -2082 347 -2048 381
rect -1964 347 -1930 381
rect -1846 347 -1812 381
rect -1728 347 -1694 381
rect -1610 347 -1576 381
rect -1492 347 -1458 381
rect -1374 347 -1340 381
rect -1256 347 -1222 381
rect -1138 347 -1104 381
rect -1020 347 -986 381
rect -902 347 -868 381
rect -784 347 -750 381
rect -666 347 -632 381
rect -548 347 -514 381
rect -430 347 -396 381
rect -312 347 -278 381
rect -194 347 -160 381
rect -76 347 -42 381
rect 42 347 76 381
rect 160 347 194 381
rect 278 347 312 381
rect 396 347 430 381
rect 514 347 548 381
rect 632 347 666 381
rect 750 347 784 381
rect 868 347 902 381
rect 986 347 1020 381
rect 1104 347 1138 381
rect 1222 347 1256 381
rect 1340 347 1374 381
rect 1458 347 1492 381
rect 1576 347 1610 381
rect 1694 347 1728 381
rect 1812 347 1846 381
rect 1930 347 1964 381
rect 2048 347 2082 381
rect 2166 347 2200 381
rect 2284 347 2318 381
rect 2402 347 2436 381
rect 2520 347 2554 381
rect 2638 347 2672 381
rect 2756 347 2790 381
rect 2874 347 2908 381
rect -2908 -381 -2874 -347
rect -2790 -381 -2756 -347
rect -2672 -381 -2638 -347
rect -2554 -381 -2520 -347
rect -2436 -381 -2402 -347
rect -2318 -381 -2284 -347
rect -2200 -381 -2166 -347
rect -2082 -381 -2048 -347
rect -1964 -381 -1930 -347
rect -1846 -381 -1812 -347
rect -1728 -381 -1694 -347
rect -1610 -381 -1576 -347
rect -1492 -381 -1458 -347
rect -1374 -381 -1340 -347
rect -1256 -381 -1222 -347
rect -1138 -381 -1104 -347
rect -1020 -381 -986 -347
rect -902 -381 -868 -347
rect -784 -381 -750 -347
rect -666 -381 -632 -347
rect -548 -381 -514 -347
rect -430 -381 -396 -347
rect -312 -381 -278 -347
rect -194 -381 -160 -347
rect -76 -381 -42 -347
rect 42 -381 76 -347
rect 160 -381 194 -347
rect 278 -381 312 -347
rect 396 -381 430 -347
rect 514 -381 548 -347
rect 632 -381 666 -347
rect 750 -381 784 -347
rect 868 -381 902 -347
rect 986 -381 1020 -347
rect 1104 -381 1138 -347
rect 1222 -381 1256 -347
rect 1340 -381 1374 -347
rect 1458 -381 1492 -347
rect 1576 -381 1610 -347
rect 1694 -381 1728 -347
rect 1812 -381 1846 -347
rect 1930 -381 1964 -347
rect 2048 -381 2082 -347
rect 2166 -381 2200 -347
rect 2284 -381 2318 -347
rect 2402 -381 2436 -347
rect 2520 -381 2554 -347
rect 2638 -381 2672 -347
rect 2756 -381 2790 -347
rect 2874 -381 2908 -347
rect -2908 -489 -2874 -455
rect -2790 -489 -2756 -455
rect -2672 -489 -2638 -455
rect -2554 -489 -2520 -455
rect -2436 -489 -2402 -455
rect -2318 -489 -2284 -455
rect -2200 -489 -2166 -455
rect -2082 -489 -2048 -455
rect -1964 -489 -1930 -455
rect -1846 -489 -1812 -455
rect -1728 -489 -1694 -455
rect -1610 -489 -1576 -455
rect -1492 -489 -1458 -455
rect -1374 -489 -1340 -455
rect -1256 -489 -1222 -455
rect -1138 -489 -1104 -455
rect -1020 -489 -986 -455
rect -902 -489 -868 -455
rect -784 -489 -750 -455
rect -666 -489 -632 -455
rect -548 -489 -514 -455
rect -430 -489 -396 -455
rect -312 -489 -278 -455
rect -194 -489 -160 -455
rect -76 -489 -42 -455
rect 42 -489 76 -455
rect 160 -489 194 -455
rect 278 -489 312 -455
rect 396 -489 430 -455
rect 514 -489 548 -455
rect 632 -489 666 -455
rect 750 -489 784 -455
rect 868 -489 902 -455
rect 986 -489 1020 -455
rect 1104 -489 1138 -455
rect 1222 -489 1256 -455
rect 1340 -489 1374 -455
rect 1458 -489 1492 -455
rect 1576 -489 1610 -455
rect 1694 -489 1728 -455
rect 1812 -489 1846 -455
rect 1930 -489 1964 -455
rect 2048 -489 2082 -455
rect 2166 -489 2200 -455
rect 2284 -489 2318 -455
rect 2402 -489 2436 -455
rect 2520 -489 2554 -455
rect 2638 -489 2672 -455
rect 2756 -489 2790 -455
rect 2874 -489 2908 -455
rect -2908 -1217 -2874 -1183
rect -2790 -1217 -2756 -1183
rect -2672 -1217 -2638 -1183
rect -2554 -1217 -2520 -1183
rect -2436 -1217 -2402 -1183
rect -2318 -1217 -2284 -1183
rect -2200 -1217 -2166 -1183
rect -2082 -1217 -2048 -1183
rect -1964 -1217 -1930 -1183
rect -1846 -1217 -1812 -1183
rect -1728 -1217 -1694 -1183
rect -1610 -1217 -1576 -1183
rect -1492 -1217 -1458 -1183
rect -1374 -1217 -1340 -1183
rect -1256 -1217 -1222 -1183
rect -1138 -1217 -1104 -1183
rect -1020 -1217 -986 -1183
rect -902 -1217 -868 -1183
rect -784 -1217 -750 -1183
rect -666 -1217 -632 -1183
rect -548 -1217 -514 -1183
rect -430 -1217 -396 -1183
rect -312 -1217 -278 -1183
rect -194 -1217 -160 -1183
rect -76 -1217 -42 -1183
rect 42 -1217 76 -1183
rect 160 -1217 194 -1183
rect 278 -1217 312 -1183
rect 396 -1217 430 -1183
rect 514 -1217 548 -1183
rect 632 -1217 666 -1183
rect 750 -1217 784 -1183
rect 868 -1217 902 -1183
rect 986 -1217 1020 -1183
rect 1104 -1217 1138 -1183
rect 1222 -1217 1256 -1183
rect 1340 -1217 1374 -1183
rect 1458 -1217 1492 -1183
rect 1576 -1217 1610 -1183
rect 1694 -1217 1728 -1183
rect 1812 -1217 1846 -1183
rect 1930 -1217 1964 -1183
rect 2048 -1217 2082 -1183
rect 2166 -1217 2200 -1183
rect 2284 -1217 2318 -1183
rect 2402 -1217 2436 -1183
rect 2520 -1217 2554 -1183
rect 2638 -1217 2672 -1183
rect 2756 -1217 2790 -1183
rect 2874 -1217 2908 -1183
<< locali >>
rect -3081 1285 -2985 1319
rect 2985 1285 3081 1319
rect -3081 1223 -3047 1285
rect 3047 1223 3081 1285
rect -2924 1183 -2908 1217
rect -2874 1183 -2858 1217
rect -2806 1183 -2790 1217
rect -2756 1183 -2740 1217
rect -2688 1183 -2672 1217
rect -2638 1183 -2622 1217
rect -2570 1183 -2554 1217
rect -2520 1183 -2504 1217
rect -2452 1183 -2436 1217
rect -2402 1183 -2386 1217
rect -2334 1183 -2318 1217
rect -2284 1183 -2268 1217
rect -2216 1183 -2200 1217
rect -2166 1183 -2150 1217
rect -2098 1183 -2082 1217
rect -2048 1183 -2032 1217
rect -1980 1183 -1964 1217
rect -1930 1183 -1914 1217
rect -1862 1183 -1846 1217
rect -1812 1183 -1796 1217
rect -1744 1183 -1728 1217
rect -1694 1183 -1678 1217
rect -1626 1183 -1610 1217
rect -1576 1183 -1560 1217
rect -1508 1183 -1492 1217
rect -1458 1183 -1442 1217
rect -1390 1183 -1374 1217
rect -1340 1183 -1324 1217
rect -1272 1183 -1256 1217
rect -1222 1183 -1206 1217
rect -1154 1183 -1138 1217
rect -1104 1183 -1088 1217
rect -1036 1183 -1020 1217
rect -986 1183 -970 1217
rect -918 1183 -902 1217
rect -868 1183 -852 1217
rect -800 1183 -784 1217
rect -750 1183 -734 1217
rect -682 1183 -666 1217
rect -632 1183 -616 1217
rect -564 1183 -548 1217
rect -514 1183 -498 1217
rect -446 1183 -430 1217
rect -396 1183 -380 1217
rect -328 1183 -312 1217
rect -278 1183 -262 1217
rect -210 1183 -194 1217
rect -160 1183 -144 1217
rect -92 1183 -76 1217
rect -42 1183 -26 1217
rect 26 1183 42 1217
rect 76 1183 92 1217
rect 144 1183 160 1217
rect 194 1183 210 1217
rect 262 1183 278 1217
rect 312 1183 328 1217
rect 380 1183 396 1217
rect 430 1183 446 1217
rect 498 1183 514 1217
rect 548 1183 564 1217
rect 616 1183 632 1217
rect 666 1183 682 1217
rect 734 1183 750 1217
rect 784 1183 800 1217
rect 852 1183 868 1217
rect 902 1183 918 1217
rect 970 1183 986 1217
rect 1020 1183 1036 1217
rect 1088 1183 1104 1217
rect 1138 1183 1154 1217
rect 1206 1183 1222 1217
rect 1256 1183 1272 1217
rect 1324 1183 1340 1217
rect 1374 1183 1390 1217
rect 1442 1183 1458 1217
rect 1492 1183 1508 1217
rect 1560 1183 1576 1217
rect 1610 1183 1626 1217
rect 1678 1183 1694 1217
rect 1728 1183 1744 1217
rect 1796 1183 1812 1217
rect 1846 1183 1862 1217
rect 1914 1183 1930 1217
rect 1964 1183 1980 1217
rect 2032 1183 2048 1217
rect 2082 1183 2098 1217
rect 2150 1183 2166 1217
rect 2200 1183 2216 1217
rect 2268 1183 2284 1217
rect 2318 1183 2334 1217
rect 2386 1183 2402 1217
rect 2436 1183 2452 1217
rect 2504 1183 2520 1217
rect 2554 1183 2570 1217
rect 2622 1183 2638 1217
rect 2672 1183 2688 1217
rect 2740 1183 2756 1217
rect 2790 1183 2806 1217
rect 2858 1183 2874 1217
rect 2908 1183 2924 1217
rect -2967 1124 -2933 1140
rect -2967 532 -2933 548
rect -2849 1124 -2815 1140
rect -2849 532 -2815 548
rect -2731 1124 -2697 1140
rect -2731 532 -2697 548
rect -2613 1124 -2579 1140
rect -2613 532 -2579 548
rect -2495 1124 -2461 1140
rect -2495 532 -2461 548
rect -2377 1124 -2343 1140
rect -2377 532 -2343 548
rect -2259 1124 -2225 1140
rect -2259 532 -2225 548
rect -2141 1124 -2107 1140
rect -2141 532 -2107 548
rect -2023 1124 -1989 1140
rect -2023 532 -1989 548
rect -1905 1124 -1871 1140
rect -1905 532 -1871 548
rect -1787 1124 -1753 1140
rect -1787 532 -1753 548
rect -1669 1124 -1635 1140
rect -1669 532 -1635 548
rect -1551 1124 -1517 1140
rect -1551 532 -1517 548
rect -1433 1124 -1399 1140
rect -1433 532 -1399 548
rect -1315 1124 -1281 1140
rect -1315 532 -1281 548
rect -1197 1124 -1163 1140
rect -1197 532 -1163 548
rect -1079 1124 -1045 1140
rect -1079 532 -1045 548
rect -961 1124 -927 1140
rect -961 532 -927 548
rect -843 1124 -809 1140
rect -843 532 -809 548
rect -725 1124 -691 1140
rect -725 532 -691 548
rect -607 1124 -573 1140
rect -607 532 -573 548
rect -489 1124 -455 1140
rect -489 532 -455 548
rect -371 1124 -337 1140
rect -371 532 -337 548
rect -253 1124 -219 1140
rect -253 532 -219 548
rect -135 1124 -101 1140
rect -135 532 -101 548
rect -17 1124 17 1140
rect -17 532 17 548
rect 101 1124 135 1140
rect 101 532 135 548
rect 219 1124 253 1140
rect 219 532 253 548
rect 337 1124 371 1140
rect 337 532 371 548
rect 455 1124 489 1140
rect 455 532 489 548
rect 573 1124 607 1140
rect 573 532 607 548
rect 691 1124 725 1140
rect 691 532 725 548
rect 809 1124 843 1140
rect 809 532 843 548
rect 927 1124 961 1140
rect 927 532 961 548
rect 1045 1124 1079 1140
rect 1045 532 1079 548
rect 1163 1124 1197 1140
rect 1163 532 1197 548
rect 1281 1124 1315 1140
rect 1281 532 1315 548
rect 1399 1124 1433 1140
rect 1399 532 1433 548
rect 1517 1124 1551 1140
rect 1517 532 1551 548
rect 1635 1124 1669 1140
rect 1635 532 1669 548
rect 1753 1124 1787 1140
rect 1753 532 1787 548
rect 1871 1124 1905 1140
rect 1871 532 1905 548
rect 1989 1124 2023 1140
rect 1989 532 2023 548
rect 2107 1124 2141 1140
rect 2107 532 2141 548
rect 2225 1124 2259 1140
rect 2225 532 2259 548
rect 2343 1124 2377 1140
rect 2343 532 2377 548
rect 2461 1124 2495 1140
rect 2461 532 2495 548
rect 2579 1124 2613 1140
rect 2579 532 2613 548
rect 2697 1124 2731 1140
rect 2697 532 2731 548
rect 2815 1124 2849 1140
rect 2815 532 2849 548
rect 2933 1124 2967 1140
rect 2933 532 2967 548
rect -2924 455 -2908 489
rect -2874 455 -2858 489
rect -2806 455 -2790 489
rect -2756 455 -2740 489
rect -2688 455 -2672 489
rect -2638 455 -2622 489
rect -2570 455 -2554 489
rect -2520 455 -2504 489
rect -2452 455 -2436 489
rect -2402 455 -2386 489
rect -2334 455 -2318 489
rect -2284 455 -2268 489
rect -2216 455 -2200 489
rect -2166 455 -2150 489
rect -2098 455 -2082 489
rect -2048 455 -2032 489
rect -1980 455 -1964 489
rect -1930 455 -1914 489
rect -1862 455 -1846 489
rect -1812 455 -1796 489
rect -1744 455 -1728 489
rect -1694 455 -1678 489
rect -1626 455 -1610 489
rect -1576 455 -1560 489
rect -1508 455 -1492 489
rect -1458 455 -1442 489
rect -1390 455 -1374 489
rect -1340 455 -1324 489
rect -1272 455 -1256 489
rect -1222 455 -1206 489
rect -1154 455 -1138 489
rect -1104 455 -1088 489
rect -1036 455 -1020 489
rect -986 455 -970 489
rect -918 455 -902 489
rect -868 455 -852 489
rect -800 455 -784 489
rect -750 455 -734 489
rect -682 455 -666 489
rect -632 455 -616 489
rect -564 455 -548 489
rect -514 455 -498 489
rect -446 455 -430 489
rect -396 455 -380 489
rect -328 455 -312 489
rect -278 455 -262 489
rect -210 455 -194 489
rect -160 455 -144 489
rect -92 455 -76 489
rect -42 455 -26 489
rect 26 455 42 489
rect 76 455 92 489
rect 144 455 160 489
rect 194 455 210 489
rect 262 455 278 489
rect 312 455 328 489
rect 380 455 396 489
rect 430 455 446 489
rect 498 455 514 489
rect 548 455 564 489
rect 616 455 632 489
rect 666 455 682 489
rect 734 455 750 489
rect 784 455 800 489
rect 852 455 868 489
rect 902 455 918 489
rect 970 455 986 489
rect 1020 455 1036 489
rect 1088 455 1104 489
rect 1138 455 1154 489
rect 1206 455 1222 489
rect 1256 455 1272 489
rect 1324 455 1340 489
rect 1374 455 1390 489
rect 1442 455 1458 489
rect 1492 455 1508 489
rect 1560 455 1576 489
rect 1610 455 1626 489
rect 1678 455 1694 489
rect 1728 455 1744 489
rect 1796 455 1812 489
rect 1846 455 1862 489
rect 1914 455 1930 489
rect 1964 455 1980 489
rect 2032 455 2048 489
rect 2082 455 2098 489
rect 2150 455 2166 489
rect 2200 455 2216 489
rect 2268 455 2284 489
rect 2318 455 2334 489
rect 2386 455 2402 489
rect 2436 455 2452 489
rect 2504 455 2520 489
rect 2554 455 2570 489
rect 2622 455 2638 489
rect 2672 455 2688 489
rect 2740 455 2756 489
rect 2790 455 2806 489
rect 2858 455 2874 489
rect 2908 455 2924 489
rect -2924 347 -2908 381
rect -2874 347 -2858 381
rect -2806 347 -2790 381
rect -2756 347 -2740 381
rect -2688 347 -2672 381
rect -2638 347 -2622 381
rect -2570 347 -2554 381
rect -2520 347 -2504 381
rect -2452 347 -2436 381
rect -2402 347 -2386 381
rect -2334 347 -2318 381
rect -2284 347 -2268 381
rect -2216 347 -2200 381
rect -2166 347 -2150 381
rect -2098 347 -2082 381
rect -2048 347 -2032 381
rect -1980 347 -1964 381
rect -1930 347 -1914 381
rect -1862 347 -1846 381
rect -1812 347 -1796 381
rect -1744 347 -1728 381
rect -1694 347 -1678 381
rect -1626 347 -1610 381
rect -1576 347 -1560 381
rect -1508 347 -1492 381
rect -1458 347 -1442 381
rect -1390 347 -1374 381
rect -1340 347 -1324 381
rect -1272 347 -1256 381
rect -1222 347 -1206 381
rect -1154 347 -1138 381
rect -1104 347 -1088 381
rect -1036 347 -1020 381
rect -986 347 -970 381
rect -918 347 -902 381
rect -868 347 -852 381
rect -800 347 -784 381
rect -750 347 -734 381
rect -682 347 -666 381
rect -632 347 -616 381
rect -564 347 -548 381
rect -514 347 -498 381
rect -446 347 -430 381
rect -396 347 -380 381
rect -328 347 -312 381
rect -278 347 -262 381
rect -210 347 -194 381
rect -160 347 -144 381
rect -92 347 -76 381
rect -42 347 -26 381
rect 26 347 42 381
rect 76 347 92 381
rect 144 347 160 381
rect 194 347 210 381
rect 262 347 278 381
rect 312 347 328 381
rect 380 347 396 381
rect 430 347 446 381
rect 498 347 514 381
rect 548 347 564 381
rect 616 347 632 381
rect 666 347 682 381
rect 734 347 750 381
rect 784 347 800 381
rect 852 347 868 381
rect 902 347 918 381
rect 970 347 986 381
rect 1020 347 1036 381
rect 1088 347 1104 381
rect 1138 347 1154 381
rect 1206 347 1222 381
rect 1256 347 1272 381
rect 1324 347 1340 381
rect 1374 347 1390 381
rect 1442 347 1458 381
rect 1492 347 1508 381
rect 1560 347 1576 381
rect 1610 347 1626 381
rect 1678 347 1694 381
rect 1728 347 1744 381
rect 1796 347 1812 381
rect 1846 347 1862 381
rect 1914 347 1930 381
rect 1964 347 1980 381
rect 2032 347 2048 381
rect 2082 347 2098 381
rect 2150 347 2166 381
rect 2200 347 2216 381
rect 2268 347 2284 381
rect 2318 347 2334 381
rect 2386 347 2402 381
rect 2436 347 2452 381
rect 2504 347 2520 381
rect 2554 347 2570 381
rect 2622 347 2638 381
rect 2672 347 2688 381
rect 2740 347 2756 381
rect 2790 347 2806 381
rect 2858 347 2874 381
rect 2908 347 2924 381
rect -2967 288 -2933 304
rect -2967 -304 -2933 -288
rect -2849 288 -2815 304
rect -2849 -304 -2815 -288
rect -2731 288 -2697 304
rect -2731 -304 -2697 -288
rect -2613 288 -2579 304
rect -2613 -304 -2579 -288
rect -2495 288 -2461 304
rect -2495 -304 -2461 -288
rect -2377 288 -2343 304
rect -2377 -304 -2343 -288
rect -2259 288 -2225 304
rect -2259 -304 -2225 -288
rect -2141 288 -2107 304
rect -2141 -304 -2107 -288
rect -2023 288 -1989 304
rect -2023 -304 -1989 -288
rect -1905 288 -1871 304
rect -1905 -304 -1871 -288
rect -1787 288 -1753 304
rect -1787 -304 -1753 -288
rect -1669 288 -1635 304
rect -1669 -304 -1635 -288
rect -1551 288 -1517 304
rect -1551 -304 -1517 -288
rect -1433 288 -1399 304
rect -1433 -304 -1399 -288
rect -1315 288 -1281 304
rect -1315 -304 -1281 -288
rect -1197 288 -1163 304
rect -1197 -304 -1163 -288
rect -1079 288 -1045 304
rect -1079 -304 -1045 -288
rect -961 288 -927 304
rect -961 -304 -927 -288
rect -843 288 -809 304
rect -843 -304 -809 -288
rect -725 288 -691 304
rect -725 -304 -691 -288
rect -607 288 -573 304
rect -607 -304 -573 -288
rect -489 288 -455 304
rect -489 -304 -455 -288
rect -371 288 -337 304
rect -371 -304 -337 -288
rect -253 288 -219 304
rect -253 -304 -219 -288
rect -135 288 -101 304
rect -135 -304 -101 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 101 288 135 304
rect 101 -304 135 -288
rect 219 288 253 304
rect 219 -304 253 -288
rect 337 288 371 304
rect 337 -304 371 -288
rect 455 288 489 304
rect 455 -304 489 -288
rect 573 288 607 304
rect 573 -304 607 -288
rect 691 288 725 304
rect 691 -304 725 -288
rect 809 288 843 304
rect 809 -304 843 -288
rect 927 288 961 304
rect 927 -304 961 -288
rect 1045 288 1079 304
rect 1045 -304 1079 -288
rect 1163 288 1197 304
rect 1163 -304 1197 -288
rect 1281 288 1315 304
rect 1281 -304 1315 -288
rect 1399 288 1433 304
rect 1399 -304 1433 -288
rect 1517 288 1551 304
rect 1517 -304 1551 -288
rect 1635 288 1669 304
rect 1635 -304 1669 -288
rect 1753 288 1787 304
rect 1753 -304 1787 -288
rect 1871 288 1905 304
rect 1871 -304 1905 -288
rect 1989 288 2023 304
rect 1989 -304 2023 -288
rect 2107 288 2141 304
rect 2107 -304 2141 -288
rect 2225 288 2259 304
rect 2225 -304 2259 -288
rect 2343 288 2377 304
rect 2343 -304 2377 -288
rect 2461 288 2495 304
rect 2461 -304 2495 -288
rect 2579 288 2613 304
rect 2579 -304 2613 -288
rect 2697 288 2731 304
rect 2697 -304 2731 -288
rect 2815 288 2849 304
rect 2815 -304 2849 -288
rect 2933 288 2967 304
rect 2933 -304 2967 -288
rect -2924 -381 -2908 -347
rect -2874 -381 -2858 -347
rect -2806 -381 -2790 -347
rect -2756 -381 -2740 -347
rect -2688 -381 -2672 -347
rect -2638 -381 -2622 -347
rect -2570 -381 -2554 -347
rect -2520 -381 -2504 -347
rect -2452 -381 -2436 -347
rect -2402 -381 -2386 -347
rect -2334 -381 -2318 -347
rect -2284 -381 -2268 -347
rect -2216 -381 -2200 -347
rect -2166 -381 -2150 -347
rect -2098 -381 -2082 -347
rect -2048 -381 -2032 -347
rect -1980 -381 -1964 -347
rect -1930 -381 -1914 -347
rect -1862 -381 -1846 -347
rect -1812 -381 -1796 -347
rect -1744 -381 -1728 -347
rect -1694 -381 -1678 -347
rect -1626 -381 -1610 -347
rect -1576 -381 -1560 -347
rect -1508 -381 -1492 -347
rect -1458 -381 -1442 -347
rect -1390 -381 -1374 -347
rect -1340 -381 -1324 -347
rect -1272 -381 -1256 -347
rect -1222 -381 -1206 -347
rect -1154 -381 -1138 -347
rect -1104 -381 -1088 -347
rect -1036 -381 -1020 -347
rect -986 -381 -970 -347
rect -918 -381 -902 -347
rect -868 -381 -852 -347
rect -800 -381 -784 -347
rect -750 -381 -734 -347
rect -682 -381 -666 -347
rect -632 -381 -616 -347
rect -564 -381 -548 -347
rect -514 -381 -498 -347
rect -446 -381 -430 -347
rect -396 -381 -380 -347
rect -328 -381 -312 -347
rect -278 -381 -262 -347
rect -210 -381 -194 -347
rect -160 -381 -144 -347
rect -92 -381 -76 -347
rect -42 -381 -26 -347
rect 26 -381 42 -347
rect 76 -381 92 -347
rect 144 -381 160 -347
rect 194 -381 210 -347
rect 262 -381 278 -347
rect 312 -381 328 -347
rect 380 -381 396 -347
rect 430 -381 446 -347
rect 498 -381 514 -347
rect 548 -381 564 -347
rect 616 -381 632 -347
rect 666 -381 682 -347
rect 734 -381 750 -347
rect 784 -381 800 -347
rect 852 -381 868 -347
rect 902 -381 918 -347
rect 970 -381 986 -347
rect 1020 -381 1036 -347
rect 1088 -381 1104 -347
rect 1138 -381 1154 -347
rect 1206 -381 1222 -347
rect 1256 -381 1272 -347
rect 1324 -381 1340 -347
rect 1374 -381 1390 -347
rect 1442 -381 1458 -347
rect 1492 -381 1508 -347
rect 1560 -381 1576 -347
rect 1610 -381 1626 -347
rect 1678 -381 1694 -347
rect 1728 -381 1744 -347
rect 1796 -381 1812 -347
rect 1846 -381 1862 -347
rect 1914 -381 1930 -347
rect 1964 -381 1980 -347
rect 2032 -381 2048 -347
rect 2082 -381 2098 -347
rect 2150 -381 2166 -347
rect 2200 -381 2216 -347
rect 2268 -381 2284 -347
rect 2318 -381 2334 -347
rect 2386 -381 2402 -347
rect 2436 -381 2452 -347
rect 2504 -381 2520 -347
rect 2554 -381 2570 -347
rect 2622 -381 2638 -347
rect 2672 -381 2688 -347
rect 2740 -381 2756 -347
rect 2790 -381 2806 -347
rect 2858 -381 2874 -347
rect 2908 -381 2924 -347
rect -2924 -489 -2908 -455
rect -2874 -489 -2858 -455
rect -2806 -489 -2790 -455
rect -2756 -489 -2740 -455
rect -2688 -489 -2672 -455
rect -2638 -489 -2622 -455
rect -2570 -489 -2554 -455
rect -2520 -489 -2504 -455
rect -2452 -489 -2436 -455
rect -2402 -489 -2386 -455
rect -2334 -489 -2318 -455
rect -2284 -489 -2268 -455
rect -2216 -489 -2200 -455
rect -2166 -489 -2150 -455
rect -2098 -489 -2082 -455
rect -2048 -489 -2032 -455
rect -1980 -489 -1964 -455
rect -1930 -489 -1914 -455
rect -1862 -489 -1846 -455
rect -1812 -489 -1796 -455
rect -1744 -489 -1728 -455
rect -1694 -489 -1678 -455
rect -1626 -489 -1610 -455
rect -1576 -489 -1560 -455
rect -1508 -489 -1492 -455
rect -1458 -489 -1442 -455
rect -1390 -489 -1374 -455
rect -1340 -489 -1324 -455
rect -1272 -489 -1256 -455
rect -1222 -489 -1206 -455
rect -1154 -489 -1138 -455
rect -1104 -489 -1088 -455
rect -1036 -489 -1020 -455
rect -986 -489 -970 -455
rect -918 -489 -902 -455
rect -868 -489 -852 -455
rect -800 -489 -784 -455
rect -750 -489 -734 -455
rect -682 -489 -666 -455
rect -632 -489 -616 -455
rect -564 -489 -548 -455
rect -514 -489 -498 -455
rect -446 -489 -430 -455
rect -396 -489 -380 -455
rect -328 -489 -312 -455
rect -278 -489 -262 -455
rect -210 -489 -194 -455
rect -160 -489 -144 -455
rect -92 -489 -76 -455
rect -42 -489 -26 -455
rect 26 -489 42 -455
rect 76 -489 92 -455
rect 144 -489 160 -455
rect 194 -489 210 -455
rect 262 -489 278 -455
rect 312 -489 328 -455
rect 380 -489 396 -455
rect 430 -489 446 -455
rect 498 -489 514 -455
rect 548 -489 564 -455
rect 616 -489 632 -455
rect 666 -489 682 -455
rect 734 -489 750 -455
rect 784 -489 800 -455
rect 852 -489 868 -455
rect 902 -489 918 -455
rect 970 -489 986 -455
rect 1020 -489 1036 -455
rect 1088 -489 1104 -455
rect 1138 -489 1154 -455
rect 1206 -489 1222 -455
rect 1256 -489 1272 -455
rect 1324 -489 1340 -455
rect 1374 -489 1390 -455
rect 1442 -489 1458 -455
rect 1492 -489 1508 -455
rect 1560 -489 1576 -455
rect 1610 -489 1626 -455
rect 1678 -489 1694 -455
rect 1728 -489 1744 -455
rect 1796 -489 1812 -455
rect 1846 -489 1862 -455
rect 1914 -489 1930 -455
rect 1964 -489 1980 -455
rect 2032 -489 2048 -455
rect 2082 -489 2098 -455
rect 2150 -489 2166 -455
rect 2200 -489 2216 -455
rect 2268 -489 2284 -455
rect 2318 -489 2334 -455
rect 2386 -489 2402 -455
rect 2436 -489 2452 -455
rect 2504 -489 2520 -455
rect 2554 -489 2570 -455
rect 2622 -489 2638 -455
rect 2672 -489 2688 -455
rect 2740 -489 2756 -455
rect 2790 -489 2806 -455
rect 2858 -489 2874 -455
rect 2908 -489 2924 -455
rect -2967 -548 -2933 -532
rect -2967 -1140 -2933 -1124
rect -2849 -548 -2815 -532
rect -2849 -1140 -2815 -1124
rect -2731 -548 -2697 -532
rect -2731 -1140 -2697 -1124
rect -2613 -548 -2579 -532
rect -2613 -1140 -2579 -1124
rect -2495 -548 -2461 -532
rect -2495 -1140 -2461 -1124
rect -2377 -548 -2343 -532
rect -2377 -1140 -2343 -1124
rect -2259 -548 -2225 -532
rect -2259 -1140 -2225 -1124
rect -2141 -548 -2107 -532
rect -2141 -1140 -2107 -1124
rect -2023 -548 -1989 -532
rect -2023 -1140 -1989 -1124
rect -1905 -548 -1871 -532
rect -1905 -1140 -1871 -1124
rect -1787 -548 -1753 -532
rect -1787 -1140 -1753 -1124
rect -1669 -548 -1635 -532
rect -1669 -1140 -1635 -1124
rect -1551 -548 -1517 -532
rect -1551 -1140 -1517 -1124
rect -1433 -548 -1399 -532
rect -1433 -1140 -1399 -1124
rect -1315 -548 -1281 -532
rect -1315 -1140 -1281 -1124
rect -1197 -548 -1163 -532
rect -1197 -1140 -1163 -1124
rect -1079 -548 -1045 -532
rect -1079 -1140 -1045 -1124
rect -961 -548 -927 -532
rect -961 -1140 -927 -1124
rect -843 -548 -809 -532
rect -843 -1140 -809 -1124
rect -725 -548 -691 -532
rect -725 -1140 -691 -1124
rect -607 -548 -573 -532
rect -607 -1140 -573 -1124
rect -489 -548 -455 -532
rect -489 -1140 -455 -1124
rect -371 -548 -337 -532
rect -371 -1140 -337 -1124
rect -253 -548 -219 -532
rect -253 -1140 -219 -1124
rect -135 -548 -101 -532
rect -135 -1140 -101 -1124
rect -17 -548 17 -532
rect -17 -1140 17 -1124
rect 101 -548 135 -532
rect 101 -1140 135 -1124
rect 219 -548 253 -532
rect 219 -1140 253 -1124
rect 337 -548 371 -532
rect 337 -1140 371 -1124
rect 455 -548 489 -532
rect 455 -1140 489 -1124
rect 573 -548 607 -532
rect 573 -1140 607 -1124
rect 691 -548 725 -532
rect 691 -1140 725 -1124
rect 809 -548 843 -532
rect 809 -1140 843 -1124
rect 927 -548 961 -532
rect 927 -1140 961 -1124
rect 1045 -548 1079 -532
rect 1045 -1140 1079 -1124
rect 1163 -548 1197 -532
rect 1163 -1140 1197 -1124
rect 1281 -548 1315 -532
rect 1281 -1140 1315 -1124
rect 1399 -548 1433 -532
rect 1399 -1140 1433 -1124
rect 1517 -548 1551 -532
rect 1517 -1140 1551 -1124
rect 1635 -548 1669 -532
rect 1635 -1140 1669 -1124
rect 1753 -548 1787 -532
rect 1753 -1140 1787 -1124
rect 1871 -548 1905 -532
rect 1871 -1140 1905 -1124
rect 1989 -548 2023 -532
rect 1989 -1140 2023 -1124
rect 2107 -548 2141 -532
rect 2107 -1140 2141 -1124
rect 2225 -548 2259 -532
rect 2225 -1140 2259 -1124
rect 2343 -548 2377 -532
rect 2343 -1140 2377 -1124
rect 2461 -548 2495 -532
rect 2461 -1140 2495 -1124
rect 2579 -548 2613 -532
rect 2579 -1140 2613 -1124
rect 2697 -548 2731 -532
rect 2697 -1140 2731 -1124
rect 2815 -548 2849 -532
rect 2815 -1140 2849 -1124
rect 2933 -548 2967 -532
rect 2933 -1140 2967 -1124
rect -2924 -1217 -2908 -1183
rect -2874 -1217 -2858 -1183
rect -2806 -1217 -2790 -1183
rect -2756 -1217 -2740 -1183
rect -2688 -1217 -2672 -1183
rect -2638 -1217 -2622 -1183
rect -2570 -1217 -2554 -1183
rect -2520 -1217 -2504 -1183
rect -2452 -1217 -2436 -1183
rect -2402 -1217 -2386 -1183
rect -2334 -1217 -2318 -1183
rect -2284 -1217 -2268 -1183
rect -2216 -1217 -2200 -1183
rect -2166 -1217 -2150 -1183
rect -2098 -1217 -2082 -1183
rect -2048 -1217 -2032 -1183
rect -1980 -1217 -1964 -1183
rect -1930 -1217 -1914 -1183
rect -1862 -1217 -1846 -1183
rect -1812 -1217 -1796 -1183
rect -1744 -1217 -1728 -1183
rect -1694 -1217 -1678 -1183
rect -1626 -1217 -1610 -1183
rect -1576 -1217 -1560 -1183
rect -1508 -1217 -1492 -1183
rect -1458 -1217 -1442 -1183
rect -1390 -1217 -1374 -1183
rect -1340 -1217 -1324 -1183
rect -1272 -1217 -1256 -1183
rect -1222 -1217 -1206 -1183
rect -1154 -1217 -1138 -1183
rect -1104 -1217 -1088 -1183
rect -1036 -1217 -1020 -1183
rect -986 -1217 -970 -1183
rect -918 -1217 -902 -1183
rect -868 -1217 -852 -1183
rect -800 -1217 -784 -1183
rect -750 -1217 -734 -1183
rect -682 -1217 -666 -1183
rect -632 -1217 -616 -1183
rect -564 -1217 -548 -1183
rect -514 -1217 -498 -1183
rect -446 -1217 -430 -1183
rect -396 -1217 -380 -1183
rect -328 -1217 -312 -1183
rect -278 -1217 -262 -1183
rect -210 -1217 -194 -1183
rect -160 -1217 -144 -1183
rect -92 -1217 -76 -1183
rect -42 -1217 -26 -1183
rect 26 -1217 42 -1183
rect 76 -1217 92 -1183
rect 144 -1217 160 -1183
rect 194 -1217 210 -1183
rect 262 -1217 278 -1183
rect 312 -1217 328 -1183
rect 380 -1217 396 -1183
rect 430 -1217 446 -1183
rect 498 -1217 514 -1183
rect 548 -1217 564 -1183
rect 616 -1217 632 -1183
rect 666 -1217 682 -1183
rect 734 -1217 750 -1183
rect 784 -1217 800 -1183
rect 852 -1217 868 -1183
rect 902 -1217 918 -1183
rect 970 -1217 986 -1183
rect 1020 -1217 1036 -1183
rect 1088 -1217 1104 -1183
rect 1138 -1217 1154 -1183
rect 1206 -1217 1222 -1183
rect 1256 -1217 1272 -1183
rect 1324 -1217 1340 -1183
rect 1374 -1217 1390 -1183
rect 1442 -1217 1458 -1183
rect 1492 -1217 1508 -1183
rect 1560 -1217 1576 -1183
rect 1610 -1217 1626 -1183
rect 1678 -1217 1694 -1183
rect 1728 -1217 1744 -1183
rect 1796 -1217 1812 -1183
rect 1846 -1217 1862 -1183
rect 1914 -1217 1930 -1183
rect 1964 -1217 1980 -1183
rect 2032 -1217 2048 -1183
rect 2082 -1217 2098 -1183
rect 2150 -1217 2166 -1183
rect 2200 -1217 2216 -1183
rect 2268 -1217 2284 -1183
rect 2318 -1217 2334 -1183
rect 2386 -1217 2402 -1183
rect 2436 -1217 2452 -1183
rect 2504 -1217 2520 -1183
rect 2554 -1217 2570 -1183
rect 2622 -1217 2638 -1183
rect 2672 -1217 2688 -1183
rect 2740 -1217 2756 -1183
rect 2790 -1217 2806 -1183
rect 2858 -1217 2874 -1183
rect 2908 -1217 2924 -1183
rect -3081 -1285 -3047 -1223
rect 3047 -1285 3081 -1223
rect -3081 -1319 -2985 -1285
rect 2985 -1319 3081 -1285
<< viali >>
rect -2908 1183 -2874 1217
rect -2790 1183 -2756 1217
rect -2672 1183 -2638 1217
rect -2554 1183 -2520 1217
rect -2436 1183 -2402 1217
rect -2318 1183 -2284 1217
rect -2200 1183 -2166 1217
rect -2082 1183 -2048 1217
rect -1964 1183 -1930 1217
rect -1846 1183 -1812 1217
rect -1728 1183 -1694 1217
rect -1610 1183 -1576 1217
rect -1492 1183 -1458 1217
rect -1374 1183 -1340 1217
rect -1256 1183 -1222 1217
rect -1138 1183 -1104 1217
rect -1020 1183 -986 1217
rect -902 1183 -868 1217
rect -784 1183 -750 1217
rect -666 1183 -632 1217
rect -548 1183 -514 1217
rect -430 1183 -396 1217
rect -312 1183 -278 1217
rect -194 1183 -160 1217
rect -76 1183 -42 1217
rect 42 1183 76 1217
rect 160 1183 194 1217
rect 278 1183 312 1217
rect 396 1183 430 1217
rect 514 1183 548 1217
rect 632 1183 666 1217
rect 750 1183 784 1217
rect 868 1183 902 1217
rect 986 1183 1020 1217
rect 1104 1183 1138 1217
rect 1222 1183 1256 1217
rect 1340 1183 1374 1217
rect 1458 1183 1492 1217
rect 1576 1183 1610 1217
rect 1694 1183 1728 1217
rect 1812 1183 1846 1217
rect 1930 1183 1964 1217
rect 2048 1183 2082 1217
rect 2166 1183 2200 1217
rect 2284 1183 2318 1217
rect 2402 1183 2436 1217
rect 2520 1183 2554 1217
rect 2638 1183 2672 1217
rect 2756 1183 2790 1217
rect 2874 1183 2908 1217
rect -2967 548 -2933 1124
rect -2849 548 -2815 1124
rect -2731 548 -2697 1124
rect -2613 548 -2579 1124
rect -2495 548 -2461 1124
rect -2377 548 -2343 1124
rect -2259 548 -2225 1124
rect -2141 548 -2107 1124
rect -2023 548 -1989 1124
rect -1905 548 -1871 1124
rect -1787 548 -1753 1124
rect -1669 548 -1635 1124
rect -1551 548 -1517 1124
rect -1433 548 -1399 1124
rect -1315 548 -1281 1124
rect -1197 548 -1163 1124
rect -1079 548 -1045 1124
rect -961 548 -927 1124
rect -843 548 -809 1124
rect -725 548 -691 1124
rect -607 548 -573 1124
rect -489 548 -455 1124
rect -371 548 -337 1124
rect -253 548 -219 1124
rect -135 548 -101 1124
rect -17 548 17 1124
rect 101 548 135 1124
rect 219 548 253 1124
rect 337 548 371 1124
rect 455 548 489 1124
rect 573 548 607 1124
rect 691 548 725 1124
rect 809 548 843 1124
rect 927 548 961 1124
rect 1045 548 1079 1124
rect 1163 548 1197 1124
rect 1281 548 1315 1124
rect 1399 548 1433 1124
rect 1517 548 1551 1124
rect 1635 548 1669 1124
rect 1753 548 1787 1124
rect 1871 548 1905 1124
rect 1989 548 2023 1124
rect 2107 548 2141 1124
rect 2225 548 2259 1124
rect 2343 548 2377 1124
rect 2461 548 2495 1124
rect 2579 548 2613 1124
rect 2697 548 2731 1124
rect 2815 548 2849 1124
rect 2933 548 2967 1124
rect -2908 455 -2874 489
rect -2790 455 -2756 489
rect -2672 455 -2638 489
rect -2554 455 -2520 489
rect -2436 455 -2402 489
rect -2318 455 -2284 489
rect -2200 455 -2166 489
rect -2082 455 -2048 489
rect -1964 455 -1930 489
rect -1846 455 -1812 489
rect -1728 455 -1694 489
rect -1610 455 -1576 489
rect -1492 455 -1458 489
rect -1374 455 -1340 489
rect -1256 455 -1222 489
rect -1138 455 -1104 489
rect -1020 455 -986 489
rect -902 455 -868 489
rect -784 455 -750 489
rect -666 455 -632 489
rect -548 455 -514 489
rect -430 455 -396 489
rect -312 455 -278 489
rect -194 455 -160 489
rect -76 455 -42 489
rect 42 455 76 489
rect 160 455 194 489
rect 278 455 312 489
rect 396 455 430 489
rect 514 455 548 489
rect 632 455 666 489
rect 750 455 784 489
rect 868 455 902 489
rect 986 455 1020 489
rect 1104 455 1138 489
rect 1222 455 1256 489
rect 1340 455 1374 489
rect 1458 455 1492 489
rect 1576 455 1610 489
rect 1694 455 1728 489
rect 1812 455 1846 489
rect 1930 455 1964 489
rect 2048 455 2082 489
rect 2166 455 2200 489
rect 2284 455 2318 489
rect 2402 455 2436 489
rect 2520 455 2554 489
rect 2638 455 2672 489
rect 2756 455 2790 489
rect 2874 455 2908 489
rect -2908 347 -2874 381
rect -2790 347 -2756 381
rect -2672 347 -2638 381
rect -2554 347 -2520 381
rect -2436 347 -2402 381
rect -2318 347 -2284 381
rect -2200 347 -2166 381
rect -2082 347 -2048 381
rect -1964 347 -1930 381
rect -1846 347 -1812 381
rect -1728 347 -1694 381
rect -1610 347 -1576 381
rect -1492 347 -1458 381
rect -1374 347 -1340 381
rect -1256 347 -1222 381
rect -1138 347 -1104 381
rect -1020 347 -986 381
rect -902 347 -868 381
rect -784 347 -750 381
rect -666 347 -632 381
rect -548 347 -514 381
rect -430 347 -396 381
rect -312 347 -278 381
rect -194 347 -160 381
rect -76 347 -42 381
rect 42 347 76 381
rect 160 347 194 381
rect 278 347 312 381
rect 396 347 430 381
rect 514 347 548 381
rect 632 347 666 381
rect 750 347 784 381
rect 868 347 902 381
rect 986 347 1020 381
rect 1104 347 1138 381
rect 1222 347 1256 381
rect 1340 347 1374 381
rect 1458 347 1492 381
rect 1576 347 1610 381
rect 1694 347 1728 381
rect 1812 347 1846 381
rect 1930 347 1964 381
rect 2048 347 2082 381
rect 2166 347 2200 381
rect 2284 347 2318 381
rect 2402 347 2436 381
rect 2520 347 2554 381
rect 2638 347 2672 381
rect 2756 347 2790 381
rect 2874 347 2908 381
rect -2967 -288 -2933 288
rect -2849 -288 -2815 288
rect -2731 -288 -2697 288
rect -2613 -288 -2579 288
rect -2495 -288 -2461 288
rect -2377 -288 -2343 288
rect -2259 -288 -2225 288
rect -2141 -288 -2107 288
rect -2023 -288 -1989 288
rect -1905 -288 -1871 288
rect -1787 -288 -1753 288
rect -1669 -288 -1635 288
rect -1551 -288 -1517 288
rect -1433 -288 -1399 288
rect -1315 -288 -1281 288
rect -1197 -288 -1163 288
rect -1079 -288 -1045 288
rect -961 -288 -927 288
rect -843 -288 -809 288
rect -725 -288 -691 288
rect -607 -288 -573 288
rect -489 -288 -455 288
rect -371 -288 -337 288
rect -253 -288 -219 288
rect -135 -288 -101 288
rect -17 -288 17 288
rect 101 -288 135 288
rect 219 -288 253 288
rect 337 -288 371 288
rect 455 -288 489 288
rect 573 -288 607 288
rect 691 -288 725 288
rect 809 -288 843 288
rect 927 -288 961 288
rect 1045 -288 1079 288
rect 1163 -288 1197 288
rect 1281 -288 1315 288
rect 1399 -288 1433 288
rect 1517 -288 1551 288
rect 1635 -288 1669 288
rect 1753 -288 1787 288
rect 1871 -288 1905 288
rect 1989 -288 2023 288
rect 2107 -288 2141 288
rect 2225 -288 2259 288
rect 2343 -288 2377 288
rect 2461 -288 2495 288
rect 2579 -288 2613 288
rect 2697 -288 2731 288
rect 2815 -288 2849 288
rect 2933 -288 2967 288
rect -2908 -381 -2874 -347
rect -2790 -381 -2756 -347
rect -2672 -381 -2638 -347
rect -2554 -381 -2520 -347
rect -2436 -381 -2402 -347
rect -2318 -381 -2284 -347
rect -2200 -381 -2166 -347
rect -2082 -381 -2048 -347
rect -1964 -381 -1930 -347
rect -1846 -381 -1812 -347
rect -1728 -381 -1694 -347
rect -1610 -381 -1576 -347
rect -1492 -381 -1458 -347
rect -1374 -381 -1340 -347
rect -1256 -381 -1222 -347
rect -1138 -381 -1104 -347
rect -1020 -381 -986 -347
rect -902 -381 -868 -347
rect -784 -381 -750 -347
rect -666 -381 -632 -347
rect -548 -381 -514 -347
rect -430 -381 -396 -347
rect -312 -381 -278 -347
rect -194 -381 -160 -347
rect -76 -381 -42 -347
rect 42 -381 76 -347
rect 160 -381 194 -347
rect 278 -381 312 -347
rect 396 -381 430 -347
rect 514 -381 548 -347
rect 632 -381 666 -347
rect 750 -381 784 -347
rect 868 -381 902 -347
rect 986 -381 1020 -347
rect 1104 -381 1138 -347
rect 1222 -381 1256 -347
rect 1340 -381 1374 -347
rect 1458 -381 1492 -347
rect 1576 -381 1610 -347
rect 1694 -381 1728 -347
rect 1812 -381 1846 -347
rect 1930 -381 1964 -347
rect 2048 -381 2082 -347
rect 2166 -381 2200 -347
rect 2284 -381 2318 -347
rect 2402 -381 2436 -347
rect 2520 -381 2554 -347
rect 2638 -381 2672 -347
rect 2756 -381 2790 -347
rect 2874 -381 2908 -347
rect -2908 -489 -2874 -455
rect -2790 -489 -2756 -455
rect -2672 -489 -2638 -455
rect -2554 -489 -2520 -455
rect -2436 -489 -2402 -455
rect -2318 -489 -2284 -455
rect -2200 -489 -2166 -455
rect -2082 -489 -2048 -455
rect -1964 -489 -1930 -455
rect -1846 -489 -1812 -455
rect -1728 -489 -1694 -455
rect -1610 -489 -1576 -455
rect -1492 -489 -1458 -455
rect -1374 -489 -1340 -455
rect -1256 -489 -1222 -455
rect -1138 -489 -1104 -455
rect -1020 -489 -986 -455
rect -902 -489 -868 -455
rect -784 -489 -750 -455
rect -666 -489 -632 -455
rect -548 -489 -514 -455
rect -430 -489 -396 -455
rect -312 -489 -278 -455
rect -194 -489 -160 -455
rect -76 -489 -42 -455
rect 42 -489 76 -455
rect 160 -489 194 -455
rect 278 -489 312 -455
rect 396 -489 430 -455
rect 514 -489 548 -455
rect 632 -489 666 -455
rect 750 -489 784 -455
rect 868 -489 902 -455
rect 986 -489 1020 -455
rect 1104 -489 1138 -455
rect 1222 -489 1256 -455
rect 1340 -489 1374 -455
rect 1458 -489 1492 -455
rect 1576 -489 1610 -455
rect 1694 -489 1728 -455
rect 1812 -489 1846 -455
rect 1930 -489 1964 -455
rect 2048 -489 2082 -455
rect 2166 -489 2200 -455
rect 2284 -489 2318 -455
rect 2402 -489 2436 -455
rect 2520 -489 2554 -455
rect 2638 -489 2672 -455
rect 2756 -489 2790 -455
rect 2874 -489 2908 -455
rect -2967 -1124 -2933 -548
rect -2849 -1124 -2815 -548
rect -2731 -1124 -2697 -548
rect -2613 -1124 -2579 -548
rect -2495 -1124 -2461 -548
rect -2377 -1124 -2343 -548
rect -2259 -1124 -2225 -548
rect -2141 -1124 -2107 -548
rect -2023 -1124 -1989 -548
rect -1905 -1124 -1871 -548
rect -1787 -1124 -1753 -548
rect -1669 -1124 -1635 -548
rect -1551 -1124 -1517 -548
rect -1433 -1124 -1399 -548
rect -1315 -1124 -1281 -548
rect -1197 -1124 -1163 -548
rect -1079 -1124 -1045 -548
rect -961 -1124 -927 -548
rect -843 -1124 -809 -548
rect -725 -1124 -691 -548
rect -607 -1124 -573 -548
rect -489 -1124 -455 -548
rect -371 -1124 -337 -548
rect -253 -1124 -219 -548
rect -135 -1124 -101 -548
rect -17 -1124 17 -548
rect 101 -1124 135 -548
rect 219 -1124 253 -548
rect 337 -1124 371 -548
rect 455 -1124 489 -548
rect 573 -1124 607 -548
rect 691 -1124 725 -548
rect 809 -1124 843 -548
rect 927 -1124 961 -548
rect 1045 -1124 1079 -548
rect 1163 -1124 1197 -548
rect 1281 -1124 1315 -548
rect 1399 -1124 1433 -548
rect 1517 -1124 1551 -548
rect 1635 -1124 1669 -548
rect 1753 -1124 1787 -548
rect 1871 -1124 1905 -548
rect 1989 -1124 2023 -548
rect 2107 -1124 2141 -548
rect 2225 -1124 2259 -548
rect 2343 -1124 2377 -548
rect 2461 -1124 2495 -548
rect 2579 -1124 2613 -548
rect 2697 -1124 2731 -548
rect 2815 -1124 2849 -548
rect 2933 -1124 2967 -548
rect -2908 -1217 -2874 -1183
rect -2790 -1217 -2756 -1183
rect -2672 -1217 -2638 -1183
rect -2554 -1217 -2520 -1183
rect -2436 -1217 -2402 -1183
rect -2318 -1217 -2284 -1183
rect -2200 -1217 -2166 -1183
rect -2082 -1217 -2048 -1183
rect -1964 -1217 -1930 -1183
rect -1846 -1217 -1812 -1183
rect -1728 -1217 -1694 -1183
rect -1610 -1217 -1576 -1183
rect -1492 -1217 -1458 -1183
rect -1374 -1217 -1340 -1183
rect -1256 -1217 -1222 -1183
rect -1138 -1217 -1104 -1183
rect -1020 -1217 -986 -1183
rect -902 -1217 -868 -1183
rect -784 -1217 -750 -1183
rect -666 -1217 -632 -1183
rect -548 -1217 -514 -1183
rect -430 -1217 -396 -1183
rect -312 -1217 -278 -1183
rect -194 -1217 -160 -1183
rect -76 -1217 -42 -1183
rect 42 -1217 76 -1183
rect 160 -1217 194 -1183
rect 278 -1217 312 -1183
rect 396 -1217 430 -1183
rect 514 -1217 548 -1183
rect 632 -1217 666 -1183
rect 750 -1217 784 -1183
rect 868 -1217 902 -1183
rect 986 -1217 1020 -1183
rect 1104 -1217 1138 -1183
rect 1222 -1217 1256 -1183
rect 1340 -1217 1374 -1183
rect 1458 -1217 1492 -1183
rect 1576 -1217 1610 -1183
rect 1694 -1217 1728 -1183
rect 1812 -1217 1846 -1183
rect 1930 -1217 1964 -1183
rect 2048 -1217 2082 -1183
rect 2166 -1217 2200 -1183
rect 2284 -1217 2318 -1183
rect 2402 -1217 2436 -1183
rect 2520 -1217 2554 -1183
rect 2638 -1217 2672 -1183
rect 2756 -1217 2790 -1183
rect 2874 -1217 2908 -1183
<< metal1 >>
rect -2920 1217 -2862 1223
rect -2920 1183 -2908 1217
rect -2874 1183 -2862 1217
rect -2920 1177 -2862 1183
rect -2802 1217 -2744 1223
rect -2802 1183 -2790 1217
rect -2756 1183 -2744 1217
rect -2802 1177 -2744 1183
rect -2684 1217 -2626 1223
rect -2684 1183 -2672 1217
rect -2638 1183 -2626 1217
rect -2684 1177 -2626 1183
rect -2566 1217 -2508 1223
rect -2566 1183 -2554 1217
rect -2520 1183 -2508 1217
rect -2566 1177 -2508 1183
rect -2448 1217 -2390 1223
rect -2448 1183 -2436 1217
rect -2402 1183 -2390 1217
rect -2448 1177 -2390 1183
rect -2330 1217 -2272 1223
rect -2330 1183 -2318 1217
rect -2284 1183 -2272 1217
rect -2330 1177 -2272 1183
rect -2212 1217 -2154 1223
rect -2212 1183 -2200 1217
rect -2166 1183 -2154 1217
rect -2212 1177 -2154 1183
rect -2094 1217 -2036 1223
rect -2094 1183 -2082 1217
rect -2048 1183 -2036 1217
rect -2094 1177 -2036 1183
rect -1976 1217 -1918 1223
rect -1976 1183 -1964 1217
rect -1930 1183 -1918 1217
rect -1976 1177 -1918 1183
rect -1858 1217 -1800 1223
rect -1858 1183 -1846 1217
rect -1812 1183 -1800 1217
rect -1858 1177 -1800 1183
rect -1740 1217 -1682 1223
rect -1740 1183 -1728 1217
rect -1694 1183 -1682 1217
rect -1740 1177 -1682 1183
rect -1622 1217 -1564 1223
rect -1622 1183 -1610 1217
rect -1576 1183 -1564 1217
rect -1622 1177 -1564 1183
rect -1504 1217 -1446 1223
rect -1504 1183 -1492 1217
rect -1458 1183 -1446 1217
rect -1504 1177 -1446 1183
rect -1386 1217 -1328 1223
rect -1386 1183 -1374 1217
rect -1340 1183 -1328 1217
rect -1386 1177 -1328 1183
rect -1268 1217 -1210 1223
rect -1268 1183 -1256 1217
rect -1222 1183 -1210 1217
rect -1268 1177 -1210 1183
rect -1150 1217 -1092 1223
rect -1150 1183 -1138 1217
rect -1104 1183 -1092 1217
rect -1150 1177 -1092 1183
rect -1032 1217 -974 1223
rect -1032 1183 -1020 1217
rect -986 1183 -974 1217
rect -1032 1177 -974 1183
rect -914 1217 -856 1223
rect -914 1183 -902 1217
rect -868 1183 -856 1217
rect -914 1177 -856 1183
rect -796 1217 -738 1223
rect -796 1183 -784 1217
rect -750 1183 -738 1217
rect -796 1177 -738 1183
rect -678 1217 -620 1223
rect -678 1183 -666 1217
rect -632 1183 -620 1217
rect -678 1177 -620 1183
rect -560 1217 -502 1223
rect -560 1183 -548 1217
rect -514 1183 -502 1217
rect -560 1177 -502 1183
rect -442 1217 -384 1223
rect -442 1183 -430 1217
rect -396 1183 -384 1217
rect -442 1177 -384 1183
rect -324 1217 -266 1223
rect -324 1183 -312 1217
rect -278 1183 -266 1217
rect -324 1177 -266 1183
rect -206 1217 -148 1223
rect -206 1183 -194 1217
rect -160 1183 -148 1217
rect -206 1177 -148 1183
rect -88 1217 -30 1223
rect -88 1183 -76 1217
rect -42 1183 -30 1217
rect -88 1177 -30 1183
rect 30 1217 88 1223
rect 30 1183 42 1217
rect 76 1183 88 1217
rect 30 1177 88 1183
rect 148 1217 206 1223
rect 148 1183 160 1217
rect 194 1183 206 1217
rect 148 1177 206 1183
rect 266 1217 324 1223
rect 266 1183 278 1217
rect 312 1183 324 1217
rect 266 1177 324 1183
rect 384 1217 442 1223
rect 384 1183 396 1217
rect 430 1183 442 1217
rect 384 1177 442 1183
rect 502 1217 560 1223
rect 502 1183 514 1217
rect 548 1183 560 1217
rect 502 1177 560 1183
rect 620 1217 678 1223
rect 620 1183 632 1217
rect 666 1183 678 1217
rect 620 1177 678 1183
rect 738 1217 796 1223
rect 738 1183 750 1217
rect 784 1183 796 1217
rect 738 1177 796 1183
rect 856 1217 914 1223
rect 856 1183 868 1217
rect 902 1183 914 1217
rect 856 1177 914 1183
rect 974 1217 1032 1223
rect 974 1183 986 1217
rect 1020 1183 1032 1217
rect 974 1177 1032 1183
rect 1092 1217 1150 1223
rect 1092 1183 1104 1217
rect 1138 1183 1150 1217
rect 1092 1177 1150 1183
rect 1210 1217 1268 1223
rect 1210 1183 1222 1217
rect 1256 1183 1268 1217
rect 1210 1177 1268 1183
rect 1328 1217 1386 1223
rect 1328 1183 1340 1217
rect 1374 1183 1386 1217
rect 1328 1177 1386 1183
rect 1446 1217 1504 1223
rect 1446 1183 1458 1217
rect 1492 1183 1504 1217
rect 1446 1177 1504 1183
rect 1564 1217 1622 1223
rect 1564 1183 1576 1217
rect 1610 1183 1622 1217
rect 1564 1177 1622 1183
rect 1682 1217 1740 1223
rect 1682 1183 1694 1217
rect 1728 1183 1740 1217
rect 1682 1177 1740 1183
rect 1800 1217 1858 1223
rect 1800 1183 1812 1217
rect 1846 1183 1858 1217
rect 1800 1177 1858 1183
rect 1918 1217 1976 1223
rect 1918 1183 1930 1217
rect 1964 1183 1976 1217
rect 1918 1177 1976 1183
rect 2036 1217 2094 1223
rect 2036 1183 2048 1217
rect 2082 1183 2094 1217
rect 2036 1177 2094 1183
rect 2154 1217 2212 1223
rect 2154 1183 2166 1217
rect 2200 1183 2212 1217
rect 2154 1177 2212 1183
rect 2272 1217 2330 1223
rect 2272 1183 2284 1217
rect 2318 1183 2330 1217
rect 2272 1177 2330 1183
rect 2390 1217 2448 1223
rect 2390 1183 2402 1217
rect 2436 1183 2448 1217
rect 2390 1177 2448 1183
rect 2508 1217 2566 1223
rect 2508 1183 2520 1217
rect 2554 1183 2566 1217
rect 2508 1177 2566 1183
rect 2626 1217 2684 1223
rect 2626 1183 2638 1217
rect 2672 1183 2684 1217
rect 2626 1177 2684 1183
rect 2744 1217 2802 1223
rect 2744 1183 2756 1217
rect 2790 1183 2802 1217
rect 2744 1177 2802 1183
rect 2862 1217 2920 1223
rect 2862 1183 2874 1217
rect 2908 1183 2920 1217
rect 2862 1177 2920 1183
rect -2973 1124 -2927 1136
rect -2973 548 -2967 1124
rect -2933 548 -2927 1124
rect -2973 536 -2927 548
rect -2855 1124 -2809 1136
rect -2855 548 -2849 1124
rect -2815 548 -2809 1124
rect -2855 536 -2809 548
rect -2737 1124 -2691 1136
rect -2737 548 -2731 1124
rect -2697 548 -2691 1124
rect -2737 536 -2691 548
rect -2619 1124 -2573 1136
rect -2619 548 -2613 1124
rect -2579 548 -2573 1124
rect -2619 536 -2573 548
rect -2501 1124 -2455 1136
rect -2501 548 -2495 1124
rect -2461 548 -2455 1124
rect -2501 536 -2455 548
rect -2383 1124 -2337 1136
rect -2383 548 -2377 1124
rect -2343 548 -2337 1124
rect -2383 536 -2337 548
rect -2265 1124 -2219 1136
rect -2265 548 -2259 1124
rect -2225 548 -2219 1124
rect -2265 536 -2219 548
rect -2147 1124 -2101 1136
rect -2147 548 -2141 1124
rect -2107 548 -2101 1124
rect -2147 536 -2101 548
rect -2029 1124 -1983 1136
rect -2029 548 -2023 1124
rect -1989 548 -1983 1124
rect -2029 536 -1983 548
rect -1911 1124 -1865 1136
rect -1911 548 -1905 1124
rect -1871 548 -1865 1124
rect -1911 536 -1865 548
rect -1793 1124 -1747 1136
rect -1793 548 -1787 1124
rect -1753 548 -1747 1124
rect -1793 536 -1747 548
rect -1675 1124 -1629 1136
rect -1675 548 -1669 1124
rect -1635 548 -1629 1124
rect -1675 536 -1629 548
rect -1557 1124 -1511 1136
rect -1557 548 -1551 1124
rect -1517 548 -1511 1124
rect -1557 536 -1511 548
rect -1439 1124 -1393 1136
rect -1439 548 -1433 1124
rect -1399 548 -1393 1124
rect -1439 536 -1393 548
rect -1321 1124 -1275 1136
rect -1321 548 -1315 1124
rect -1281 548 -1275 1124
rect -1321 536 -1275 548
rect -1203 1124 -1157 1136
rect -1203 548 -1197 1124
rect -1163 548 -1157 1124
rect -1203 536 -1157 548
rect -1085 1124 -1039 1136
rect -1085 548 -1079 1124
rect -1045 548 -1039 1124
rect -1085 536 -1039 548
rect -967 1124 -921 1136
rect -967 548 -961 1124
rect -927 548 -921 1124
rect -967 536 -921 548
rect -849 1124 -803 1136
rect -849 548 -843 1124
rect -809 548 -803 1124
rect -849 536 -803 548
rect -731 1124 -685 1136
rect -731 548 -725 1124
rect -691 548 -685 1124
rect -731 536 -685 548
rect -613 1124 -567 1136
rect -613 548 -607 1124
rect -573 548 -567 1124
rect -613 536 -567 548
rect -495 1124 -449 1136
rect -495 548 -489 1124
rect -455 548 -449 1124
rect -495 536 -449 548
rect -377 1124 -331 1136
rect -377 548 -371 1124
rect -337 548 -331 1124
rect -377 536 -331 548
rect -259 1124 -213 1136
rect -259 548 -253 1124
rect -219 548 -213 1124
rect -259 536 -213 548
rect -141 1124 -95 1136
rect -141 548 -135 1124
rect -101 548 -95 1124
rect -141 536 -95 548
rect -23 1124 23 1136
rect -23 548 -17 1124
rect 17 548 23 1124
rect -23 536 23 548
rect 95 1124 141 1136
rect 95 548 101 1124
rect 135 548 141 1124
rect 95 536 141 548
rect 213 1124 259 1136
rect 213 548 219 1124
rect 253 548 259 1124
rect 213 536 259 548
rect 331 1124 377 1136
rect 331 548 337 1124
rect 371 548 377 1124
rect 331 536 377 548
rect 449 1124 495 1136
rect 449 548 455 1124
rect 489 548 495 1124
rect 449 536 495 548
rect 567 1124 613 1136
rect 567 548 573 1124
rect 607 548 613 1124
rect 567 536 613 548
rect 685 1124 731 1136
rect 685 548 691 1124
rect 725 548 731 1124
rect 685 536 731 548
rect 803 1124 849 1136
rect 803 548 809 1124
rect 843 548 849 1124
rect 803 536 849 548
rect 921 1124 967 1136
rect 921 548 927 1124
rect 961 548 967 1124
rect 921 536 967 548
rect 1039 1124 1085 1136
rect 1039 548 1045 1124
rect 1079 548 1085 1124
rect 1039 536 1085 548
rect 1157 1124 1203 1136
rect 1157 548 1163 1124
rect 1197 548 1203 1124
rect 1157 536 1203 548
rect 1275 1124 1321 1136
rect 1275 548 1281 1124
rect 1315 548 1321 1124
rect 1275 536 1321 548
rect 1393 1124 1439 1136
rect 1393 548 1399 1124
rect 1433 548 1439 1124
rect 1393 536 1439 548
rect 1511 1124 1557 1136
rect 1511 548 1517 1124
rect 1551 548 1557 1124
rect 1511 536 1557 548
rect 1629 1124 1675 1136
rect 1629 548 1635 1124
rect 1669 548 1675 1124
rect 1629 536 1675 548
rect 1747 1124 1793 1136
rect 1747 548 1753 1124
rect 1787 548 1793 1124
rect 1747 536 1793 548
rect 1865 1124 1911 1136
rect 1865 548 1871 1124
rect 1905 548 1911 1124
rect 1865 536 1911 548
rect 1983 1124 2029 1136
rect 1983 548 1989 1124
rect 2023 548 2029 1124
rect 1983 536 2029 548
rect 2101 1124 2147 1136
rect 2101 548 2107 1124
rect 2141 548 2147 1124
rect 2101 536 2147 548
rect 2219 1124 2265 1136
rect 2219 548 2225 1124
rect 2259 548 2265 1124
rect 2219 536 2265 548
rect 2337 1124 2383 1136
rect 2337 548 2343 1124
rect 2377 548 2383 1124
rect 2337 536 2383 548
rect 2455 1124 2501 1136
rect 2455 548 2461 1124
rect 2495 548 2501 1124
rect 2455 536 2501 548
rect 2573 1124 2619 1136
rect 2573 548 2579 1124
rect 2613 548 2619 1124
rect 2573 536 2619 548
rect 2691 1124 2737 1136
rect 2691 548 2697 1124
rect 2731 548 2737 1124
rect 2691 536 2737 548
rect 2809 1124 2855 1136
rect 2809 548 2815 1124
rect 2849 548 2855 1124
rect 2809 536 2855 548
rect 2927 1124 2973 1136
rect 2927 548 2933 1124
rect 2967 548 2973 1124
rect 2927 536 2973 548
rect -2920 489 -2862 495
rect -2920 455 -2908 489
rect -2874 455 -2862 489
rect -2920 449 -2862 455
rect -2802 489 -2744 495
rect -2802 455 -2790 489
rect -2756 455 -2744 489
rect -2802 449 -2744 455
rect -2684 489 -2626 495
rect -2684 455 -2672 489
rect -2638 455 -2626 489
rect -2684 449 -2626 455
rect -2566 489 -2508 495
rect -2566 455 -2554 489
rect -2520 455 -2508 489
rect -2566 449 -2508 455
rect -2448 489 -2390 495
rect -2448 455 -2436 489
rect -2402 455 -2390 489
rect -2448 449 -2390 455
rect -2330 489 -2272 495
rect -2330 455 -2318 489
rect -2284 455 -2272 489
rect -2330 449 -2272 455
rect -2212 489 -2154 495
rect -2212 455 -2200 489
rect -2166 455 -2154 489
rect -2212 449 -2154 455
rect -2094 489 -2036 495
rect -2094 455 -2082 489
rect -2048 455 -2036 489
rect -2094 449 -2036 455
rect -1976 489 -1918 495
rect -1976 455 -1964 489
rect -1930 455 -1918 489
rect -1976 449 -1918 455
rect -1858 489 -1800 495
rect -1858 455 -1846 489
rect -1812 455 -1800 489
rect -1858 449 -1800 455
rect -1740 489 -1682 495
rect -1740 455 -1728 489
rect -1694 455 -1682 489
rect -1740 449 -1682 455
rect -1622 489 -1564 495
rect -1622 455 -1610 489
rect -1576 455 -1564 489
rect -1622 449 -1564 455
rect -1504 489 -1446 495
rect -1504 455 -1492 489
rect -1458 455 -1446 489
rect -1504 449 -1446 455
rect -1386 489 -1328 495
rect -1386 455 -1374 489
rect -1340 455 -1328 489
rect -1386 449 -1328 455
rect -1268 489 -1210 495
rect -1268 455 -1256 489
rect -1222 455 -1210 489
rect -1268 449 -1210 455
rect -1150 489 -1092 495
rect -1150 455 -1138 489
rect -1104 455 -1092 489
rect -1150 449 -1092 455
rect -1032 489 -974 495
rect -1032 455 -1020 489
rect -986 455 -974 489
rect -1032 449 -974 455
rect -914 489 -856 495
rect -914 455 -902 489
rect -868 455 -856 489
rect -914 449 -856 455
rect -796 489 -738 495
rect -796 455 -784 489
rect -750 455 -738 489
rect -796 449 -738 455
rect -678 489 -620 495
rect -678 455 -666 489
rect -632 455 -620 489
rect -678 449 -620 455
rect -560 489 -502 495
rect -560 455 -548 489
rect -514 455 -502 489
rect -560 449 -502 455
rect -442 489 -384 495
rect -442 455 -430 489
rect -396 455 -384 489
rect -442 449 -384 455
rect -324 489 -266 495
rect -324 455 -312 489
rect -278 455 -266 489
rect -324 449 -266 455
rect -206 489 -148 495
rect -206 455 -194 489
rect -160 455 -148 489
rect -206 449 -148 455
rect -88 489 -30 495
rect -88 455 -76 489
rect -42 455 -30 489
rect -88 449 -30 455
rect 30 489 88 495
rect 30 455 42 489
rect 76 455 88 489
rect 30 449 88 455
rect 148 489 206 495
rect 148 455 160 489
rect 194 455 206 489
rect 148 449 206 455
rect 266 489 324 495
rect 266 455 278 489
rect 312 455 324 489
rect 266 449 324 455
rect 384 489 442 495
rect 384 455 396 489
rect 430 455 442 489
rect 384 449 442 455
rect 502 489 560 495
rect 502 455 514 489
rect 548 455 560 489
rect 502 449 560 455
rect 620 489 678 495
rect 620 455 632 489
rect 666 455 678 489
rect 620 449 678 455
rect 738 489 796 495
rect 738 455 750 489
rect 784 455 796 489
rect 738 449 796 455
rect 856 489 914 495
rect 856 455 868 489
rect 902 455 914 489
rect 856 449 914 455
rect 974 489 1032 495
rect 974 455 986 489
rect 1020 455 1032 489
rect 974 449 1032 455
rect 1092 489 1150 495
rect 1092 455 1104 489
rect 1138 455 1150 489
rect 1092 449 1150 455
rect 1210 489 1268 495
rect 1210 455 1222 489
rect 1256 455 1268 489
rect 1210 449 1268 455
rect 1328 489 1386 495
rect 1328 455 1340 489
rect 1374 455 1386 489
rect 1328 449 1386 455
rect 1446 489 1504 495
rect 1446 455 1458 489
rect 1492 455 1504 489
rect 1446 449 1504 455
rect 1564 489 1622 495
rect 1564 455 1576 489
rect 1610 455 1622 489
rect 1564 449 1622 455
rect 1682 489 1740 495
rect 1682 455 1694 489
rect 1728 455 1740 489
rect 1682 449 1740 455
rect 1800 489 1858 495
rect 1800 455 1812 489
rect 1846 455 1858 489
rect 1800 449 1858 455
rect 1918 489 1976 495
rect 1918 455 1930 489
rect 1964 455 1976 489
rect 1918 449 1976 455
rect 2036 489 2094 495
rect 2036 455 2048 489
rect 2082 455 2094 489
rect 2036 449 2094 455
rect 2154 489 2212 495
rect 2154 455 2166 489
rect 2200 455 2212 489
rect 2154 449 2212 455
rect 2272 489 2330 495
rect 2272 455 2284 489
rect 2318 455 2330 489
rect 2272 449 2330 455
rect 2390 489 2448 495
rect 2390 455 2402 489
rect 2436 455 2448 489
rect 2390 449 2448 455
rect 2508 489 2566 495
rect 2508 455 2520 489
rect 2554 455 2566 489
rect 2508 449 2566 455
rect 2626 489 2684 495
rect 2626 455 2638 489
rect 2672 455 2684 489
rect 2626 449 2684 455
rect 2744 489 2802 495
rect 2744 455 2756 489
rect 2790 455 2802 489
rect 2744 449 2802 455
rect 2862 489 2920 495
rect 2862 455 2874 489
rect 2908 455 2920 489
rect 2862 449 2920 455
rect -2920 381 -2862 387
rect -2920 347 -2908 381
rect -2874 347 -2862 381
rect -2920 341 -2862 347
rect -2802 381 -2744 387
rect -2802 347 -2790 381
rect -2756 347 -2744 381
rect -2802 341 -2744 347
rect -2684 381 -2626 387
rect -2684 347 -2672 381
rect -2638 347 -2626 381
rect -2684 341 -2626 347
rect -2566 381 -2508 387
rect -2566 347 -2554 381
rect -2520 347 -2508 381
rect -2566 341 -2508 347
rect -2448 381 -2390 387
rect -2448 347 -2436 381
rect -2402 347 -2390 381
rect -2448 341 -2390 347
rect -2330 381 -2272 387
rect -2330 347 -2318 381
rect -2284 347 -2272 381
rect -2330 341 -2272 347
rect -2212 381 -2154 387
rect -2212 347 -2200 381
rect -2166 347 -2154 381
rect -2212 341 -2154 347
rect -2094 381 -2036 387
rect -2094 347 -2082 381
rect -2048 347 -2036 381
rect -2094 341 -2036 347
rect -1976 381 -1918 387
rect -1976 347 -1964 381
rect -1930 347 -1918 381
rect -1976 341 -1918 347
rect -1858 381 -1800 387
rect -1858 347 -1846 381
rect -1812 347 -1800 381
rect -1858 341 -1800 347
rect -1740 381 -1682 387
rect -1740 347 -1728 381
rect -1694 347 -1682 381
rect -1740 341 -1682 347
rect -1622 381 -1564 387
rect -1622 347 -1610 381
rect -1576 347 -1564 381
rect -1622 341 -1564 347
rect -1504 381 -1446 387
rect -1504 347 -1492 381
rect -1458 347 -1446 381
rect -1504 341 -1446 347
rect -1386 381 -1328 387
rect -1386 347 -1374 381
rect -1340 347 -1328 381
rect -1386 341 -1328 347
rect -1268 381 -1210 387
rect -1268 347 -1256 381
rect -1222 347 -1210 381
rect -1268 341 -1210 347
rect -1150 381 -1092 387
rect -1150 347 -1138 381
rect -1104 347 -1092 381
rect -1150 341 -1092 347
rect -1032 381 -974 387
rect -1032 347 -1020 381
rect -986 347 -974 381
rect -1032 341 -974 347
rect -914 381 -856 387
rect -914 347 -902 381
rect -868 347 -856 381
rect -914 341 -856 347
rect -796 381 -738 387
rect -796 347 -784 381
rect -750 347 -738 381
rect -796 341 -738 347
rect -678 381 -620 387
rect -678 347 -666 381
rect -632 347 -620 381
rect -678 341 -620 347
rect -560 381 -502 387
rect -560 347 -548 381
rect -514 347 -502 381
rect -560 341 -502 347
rect -442 381 -384 387
rect -442 347 -430 381
rect -396 347 -384 381
rect -442 341 -384 347
rect -324 381 -266 387
rect -324 347 -312 381
rect -278 347 -266 381
rect -324 341 -266 347
rect -206 381 -148 387
rect -206 347 -194 381
rect -160 347 -148 381
rect -206 341 -148 347
rect -88 381 -30 387
rect -88 347 -76 381
rect -42 347 -30 381
rect -88 341 -30 347
rect 30 381 88 387
rect 30 347 42 381
rect 76 347 88 381
rect 30 341 88 347
rect 148 381 206 387
rect 148 347 160 381
rect 194 347 206 381
rect 148 341 206 347
rect 266 381 324 387
rect 266 347 278 381
rect 312 347 324 381
rect 266 341 324 347
rect 384 381 442 387
rect 384 347 396 381
rect 430 347 442 381
rect 384 341 442 347
rect 502 381 560 387
rect 502 347 514 381
rect 548 347 560 381
rect 502 341 560 347
rect 620 381 678 387
rect 620 347 632 381
rect 666 347 678 381
rect 620 341 678 347
rect 738 381 796 387
rect 738 347 750 381
rect 784 347 796 381
rect 738 341 796 347
rect 856 381 914 387
rect 856 347 868 381
rect 902 347 914 381
rect 856 341 914 347
rect 974 381 1032 387
rect 974 347 986 381
rect 1020 347 1032 381
rect 974 341 1032 347
rect 1092 381 1150 387
rect 1092 347 1104 381
rect 1138 347 1150 381
rect 1092 341 1150 347
rect 1210 381 1268 387
rect 1210 347 1222 381
rect 1256 347 1268 381
rect 1210 341 1268 347
rect 1328 381 1386 387
rect 1328 347 1340 381
rect 1374 347 1386 381
rect 1328 341 1386 347
rect 1446 381 1504 387
rect 1446 347 1458 381
rect 1492 347 1504 381
rect 1446 341 1504 347
rect 1564 381 1622 387
rect 1564 347 1576 381
rect 1610 347 1622 381
rect 1564 341 1622 347
rect 1682 381 1740 387
rect 1682 347 1694 381
rect 1728 347 1740 381
rect 1682 341 1740 347
rect 1800 381 1858 387
rect 1800 347 1812 381
rect 1846 347 1858 381
rect 1800 341 1858 347
rect 1918 381 1976 387
rect 1918 347 1930 381
rect 1964 347 1976 381
rect 1918 341 1976 347
rect 2036 381 2094 387
rect 2036 347 2048 381
rect 2082 347 2094 381
rect 2036 341 2094 347
rect 2154 381 2212 387
rect 2154 347 2166 381
rect 2200 347 2212 381
rect 2154 341 2212 347
rect 2272 381 2330 387
rect 2272 347 2284 381
rect 2318 347 2330 381
rect 2272 341 2330 347
rect 2390 381 2448 387
rect 2390 347 2402 381
rect 2436 347 2448 381
rect 2390 341 2448 347
rect 2508 381 2566 387
rect 2508 347 2520 381
rect 2554 347 2566 381
rect 2508 341 2566 347
rect 2626 381 2684 387
rect 2626 347 2638 381
rect 2672 347 2684 381
rect 2626 341 2684 347
rect 2744 381 2802 387
rect 2744 347 2756 381
rect 2790 347 2802 381
rect 2744 341 2802 347
rect 2862 381 2920 387
rect 2862 347 2874 381
rect 2908 347 2920 381
rect 2862 341 2920 347
rect -2973 288 -2927 300
rect -2973 -288 -2967 288
rect -2933 -288 -2927 288
rect -2973 -300 -2927 -288
rect -2855 288 -2809 300
rect -2855 -288 -2849 288
rect -2815 -288 -2809 288
rect -2855 -300 -2809 -288
rect -2737 288 -2691 300
rect -2737 -288 -2731 288
rect -2697 -288 -2691 288
rect -2737 -300 -2691 -288
rect -2619 288 -2573 300
rect -2619 -288 -2613 288
rect -2579 -288 -2573 288
rect -2619 -300 -2573 -288
rect -2501 288 -2455 300
rect -2501 -288 -2495 288
rect -2461 -288 -2455 288
rect -2501 -300 -2455 -288
rect -2383 288 -2337 300
rect -2383 -288 -2377 288
rect -2343 -288 -2337 288
rect -2383 -300 -2337 -288
rect -2265 288 -2219 300
rect -2265 -288 -2259 288
rect -2225 -288 -2219 288
rect -2265 -300 -2219 -288
rect -2147 288 -2101 300
rect -2147 -288 -2141 288
rect -2107 -288 -2101 288
rect -2147 -300 -2101 -288
rect -2029 288 -1983 300
rect -2029 -288 -2023 288
rect -1989 -288 -1983 288
rect -2029 -300 -1983 -288
rect -1911 288 -1865 300
rect -1911 -288 -1905 288
rect -1871 -288 -1865 288
rect -1911 -300 -1865 -288
rect -1793 288 -1747 300
rect -1793 -288 -1787 288
rect -1753 -288 -1747 288
rect -1793 -300 -1747 -288
rect -1675 288 -1629 300
rect -1675 -288 -1669 288
rect -1635 -288 -1629 288
rect -1675 -300 -1629 -288
rect -1557 288 -1511 300
rect -1557 -288 -1551 288
rect -1517 -288 -1511 288
rect -1557 -300 -1511 -288
rect -1439 288 -1393 300
rect -1439 -288 -1433 288
rect -1399 -288 -1393 288
rect -1439 -300 -1393 -288
rect -1321 288 -1275 300
rect -1321 -288 -1315 288
rect -1281 -288 -1275 288
rect -1321 -300 -1275 -288
rect -1203 288 -1157 300
rect -1203 -288 -1197 288
rect -1163 -288 -1157 288
rect -1203 -300 -1157 -288
rect -1085 288 -1039 300
rect -1085 -288 -1079 288
rect -1045 -288 -1039 288
rect -1085 -300 -1039 -288
rect -967 288 -921 300
rect -967 -288 -961 288
rect -927 -288 -921 288
rect -967 -300 -921 -288
rect -849 288 -803 300
rect -849 -288 -843 288
rect -809 -288 -803 288
rect -849 -300 -803 -288
rect -731 288 -685 300
rect -731 -288 -725 288
rect -691 -288 -685 288
rect -731 -300 -685 -288
rect -613 288 -567 300
rect -613 -288 -607 288
rect -573 -288 -567 288
rect -613 -300 -567 -288
rect -495 288 -449 300
rect -495 -288 -489 288
rect -455 -288 -449 288
rect -495 -300 -449 -288
rect -377 288 -331 300
rect -377 -288 -371 288
rect -337 -288 -331 288
rect -377 -300 -331 -288
rect -259 288 -213 300
rect -259 -288 -253 288
rect -219 -288 -213 288
rect -259 -300 -213 -288
rect -141 288 -95 300
rect -141 -288 -135 288
rect -101 -288 -95 288
rect -141 -300 -95 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 95 288 141 300
rect 95 -288 101 288
rect 135 -288 141 288
rect 95 -300 141 -288
rect 213 288 259 300
rect 213 -288 219 288
rect 253 -288 259 288
rect 213 -300 259 -288
rect 331 288 377 300
rect 331 -288 337 288
rect 371 -288 377 288
rect 331 -300 377 -288
rect 449 288 495 300
rect 449 -288 455 288
rect 489 -288 495 288
rect 449 -300 495 -288
rect 567 288 613 300
rect 567 -288 573 288
rect 607 -288 613 288
rect 567 -300 613 -288
rect 685 288 731 300
rect 685 -288 691 288
rect 725 -288 731 288
rect 685 -300 731 -288
rect 803 288 849 300
rect 803 -288 809 288
rect 843 -288 849 288
rect 803 -300 849 -288
rect 921 288 967 300
rect 921 -288 927 288
rect 961 -288 967 288
rect 921 -300 967 -288
rect 1039 288 1085 300
rect 1039 -288 1045 288
rect 1079 -288 1085 288
rect 1039 -300 1085 -288
rect 1157 288 1203 300
rect 1157 -288 1163 288
rect 1197 -288 1203 288
rect 1157 -300 1203 -288
rect 1275 288 1321 300
rect 1275 -288 1281 288
rect 1315 -288 1321 288
rect 1275 -300 1321 -288
rect 1393 288 1439 300
rect 1393 -288 1399 288
rect 1433 -288 1439 288
rect 1393 -300 1439 -288
rect 1511 288 1557 300
rect 1511 -288 1517 288
rect 1551 -288 1557 288
rect 1511 -300 1557 -288
rect 1629 288 1675 300
rect 1629 -288 1635 288
rect 1669 -288 1675 288
rect 1629 -300 1675 -288
rect 1747 288 1793 300
rect 1747 -288 1753 288
rect 1787 -288 1793 288
rect 1747 -300 1793 -288
rect 1865 288 1911 300
rect 1865 -288 1871 288
rect 1905 -288 1911 288
rect 1865 -300 1911 -288
rect 1983 288 2029 300
rect 1983 -288 1989 288
rect 2023 -288 2029 288
rect 1983 -300 2029 -288
rect 2101 288 2147 300
rect 2101 -288 2107 288
rect 2141 -288 2147 288
rect 2101 -300 2147 -288
rect 2219 288 2265 300
rect 2219 -288 2225 288
rect 2259 -288 2265 288
rect 2219 -300 2265 -288
rect 2337 288 2383 300
rect 2337 -288 2343 288
rect 2377 -288 2383 288
rect 2337 -300 2383 -288
rect 2455 288 2501 300
rect 2455 -288 2461 288
rect 2495 -288 2501 288
rect 2455 -300 2501 -288
rect 2573 288 2619 300
rect 2573 -288 2579 288
rect 2613 -288 2619 288
rect 2573 -300 2619 -288
rect 2691 288 2737 300
rect 2691 -288 2697 288
rect 2731 -288 2737 288
rect 2691 -300 2737 -288
rect 2809 288 2855 300
rect 2809 -288 2815 288
rect 2849 -288 2855 288
rect 2809 -300 2855 -288
rect 2927 288 2973 300
rect 2927 -288 2933 288
rect 2967 -288 2973 288
rect 2927 -300 2973 -288
rect -2920 -347 -2862 -341
rect -2920 -381 -2908 -347
rect -2874 -381 -2862 -347
rect -2920 -387 -2862 -381
rect -2802 -347 -2744 -341
rect -2802 -381 -2790 -347
rect -2756 -381 -2744 -347
rect -2802 -387 -2744 -381
rect -2684 -347 -2626 -341
rect -2684 -381 -2672 -347
rect -2638 -381 -2626 -347
rect -2684 -387 -2626 -381
rect -2566 -347 -2508 -341
rect -2566 -381 -2554 -347
rect -2520 -381 -2508 -347
rect -2566 -387 -2508 -381
rect -2448 -347 -2390 -341
rect -2448 -381 -2436 -347
rect -2402 -381 -2390 -347
rect -2448 -387 -2390 -381
rect -2330 -347 -2272 -341
rect -2330 -381 -2318 -347
rect -2284 -381 -2272 -347
rect -2330 -387 -2272 -381
rect -2212 -347 -2154 -341
rect -2212 -381 -2200 -347
rect -2166 -381 -2154 -347
rect -2212 -387 -2154 -381
rect -2094 -347 -2036 -341
rect -2094 -381 -2082 -347
rect -2048 -381 -2036 -347
rect -2094 -387 -2036 -381
rect -1976 -347 -1918 -341
rect -1976 -381 -1964 -347
rect -1930 -381 -1918 -347
rect -1976 -387 -1918 -381
rect -1858 -347 -1800 -341
rect -1858 -381 -1846 -347
rect -1812 -381 -1800 -347
rect -1858 -387 -1800 -381
rect -1740 -347 -1682 -341
rect -1740 -381 -1728 -347
rect -1694 -381 -1682 -347
rect -1740 -387 -1682 -381
rect -1622 -347 -1564 -341
rect -1622 -381 -1610 -347
rect -1576 -381 -1564 -347
rect -1622 -387 -1564 -381
rect -1504 -347 -1446 -341
rect -1504 -381 -1492 -347
rect -1458 -381 -1446 -347
rect -1504 -387 -1446 -381
rect -1386 -347 -1328 -341
rect -1386 -381 -1374 -347
rect -1340 -381 -1328 -347
rect -1386 -387 -1328 -381
rect -1268 -347 -1210 -341
rect -1268 -381 -1256 -347
rect -1222 -381 -1210 -347
rect -1268 -387 -1210 -381
rect -1150 -347 -1092 -341
rect -1150 -381 -1138 -347
rect -1104 -381 -1092 -347
rect -1150 -387 -1092 -381
rect -1032 -347 -974 -341
rect -1032 -381 -1020 -347
rect -986 -381 -974 -347
rect -1032 -387 -974 -381
rect -914 -347 -856 -341
rect -914 -381 -902 -347
rect -868 -381 -856 -347
rect -914 -387 -856 -381
rect -796 -347 -738 -341
rect -796 -381 -784 -347
rect -750 -381 -738 -347
rect -796 -387 -738 -381
rect -678 -347 -620 -341
rect -678 -381 -666 -347
rect -632 -381 -620 -347
rect -678 -387 -620 -381
rect -560 -347 -502 -341
rect -560 -381 -548 -347
rect -514 -381 -502 -347
rect -560 -387 -502 -381
rect -442 -347 -384 -341
rect -442 -381 -430 -347
rect -396 -381 -384 -347
rect -442 -387 -384 -381
rect -324 -347 -266 -341
rect -324 -381 -312 -347
rect -278 -381 -266 -347
rect -324 -387 -266 -381
rect -206 -347 -148 -341
rect -206 -381 -194 -347
rect -160 -381 -148 -347
rect -206 -387 -148 -381
rect -88 -347 -30 -341
rect -88 -381 -76 -347
rect -42 -381 -30 -347
rect -88 -387 -30 -381
rect 30 -347 88 -341
rect 30 -381 42 -347
rect 76 -381 88 -347
rect 30 -387 88 -381
rect 148 -347 206 -341
rect 148 -381 160 -347
rect 194 -381 206 -347
rect 148 -387 206 -381
rect 266 -347 324 -341
rect 266 -381 278 -347
rect 312 -381 324 -347
rect 266 -387 324 -381
rect 384 -347 442 -341
rect 384 -381 396 -347
rect 430 -381 442 -347
rect 384 -387 442 -381
rect 502 -347 560 -341
rect 502 -381 514 -347
rect 548 -381 560 -347
rect 502 -387 560 -381
rect 620 -347 678 -341
rect 620 -381 632 -347
rect 666 -381 678 -347
rect 620 -387 678 -381
rect 738 -347 796 -341
rect 738 -381 750 -347
rect 784 -381 796 -347
rect 738 -387 796 -381
rect 856 -347 914 -341
rect 856 -381 868 -347
rect 902 -381 914 -347
rect 856 -387 914 -381
rect 974 -347 1032 -341
rect 974 -381 986 -347
rect 1020 -381 1032 -347
rect 974 -387 1032 -381
rect 1092 -347 1150 -341
rect 1092 -381 1104 -347
rect 1138 -381 1150 -347
rect 1092 -387 1150 -381
rect 1210 -347 1268 -341
rect 1210 -381 1222 -347
rect 1256 -381 1268 -347
rect 1210 -387 1268 -381
rect 1328 -347 1386 -341
rect 1328 -381 1340 -347
rect 1374 -381 1386 -347
rect 1328 -387 1386 -381
rect 1446 -347 1504 -341
rect 1446 -381 1458 -347
rect 1492 -381 1504 -347
rect 1446 -387 1504 -381
rect 1564 -347 1622 -341
rect 1564 -381 1576 -347
rect 1610 -381 1622 -347
rect 1564 -387 1622 -381
rect 1682 -347 1740 -341
rect 1682 -381 1694 -347
rect 1728 -381 1740 -347
rect 1682 -387 1740 -381
rect 1800 -347 1858 -341
rect 1800 -381 1812 -347
rect 1846 -381 1858 -347
rect 1800 -387 1858 -381
rect 1918 -347 1976 -341
rect 1918 -381 1930 -347
rect 1964 -381 1976 -347
rect 1918 -387 1976 -381
rect 2036 -347 2094 -341
rect 2036 -381 2048 -347
rect 2082 -381 2094 -347
rect 2036 -387 2094 -381
rect 2154 -347 2212 -341
rect 2154 -381 2166 -347
rect 2200 -381 2212 -347
rect 2154 -387 2212 -381
rect 2272 -347 2330 -341
rect 2272 -381 2284 -347
rect 2318 -381 2330 -347
rect 2272 -387 2330 -381
rect 2390 -347 2448 -341
rect 2390 -381 2402 -347
rect 2436 -381 2448 -347
rect 2390 -387 2448 -381
rect 2508 -347 2566 -341
rect 2508 -381 2520 -347
rect 2554 -381 2566 -347
rect 2508 -387 2566 -381
rect 2626 -347 2684 -341
rect 2626 -381 2638 -347
rect 2672 -381 2684 -347
rect 2626 -387 2684 -381
rect 2744 -347 2802 -341
rect 2744 -381 2756 -347
rect 2790 -381 2802 -347
rect 2744 -387 2802 -381
rect 2862 -347 2920 -341
rect 2862 -381 2874 -347
rect 2908 -381 2920 -347
rect 2862 -387 2920 -381
rect -2920 -455 -2862 -449
rect -2920 -489 -2908 -455
rect -2874 -489 -2862 -455
rect -2920 -495 -2862 -489
rect -2802 -455 -2744 -449
rect -2802 -489 -2790 -455
rect -2756 -489 -2744 -455
rect -2802 -495 -2744 -489
rect -2684 -455 -2626 -449
rect -2684 -489 -2672 -455
rect -2638 -489 -2626 -455
rect -2684 -495 -2626 -489
rect -2566 -455 -2508 -449
rect -2566 -489 -2554 -455
rect -2520 -489 -2508 -455
rect -2566 -495 -2508 -489
rect -2448 -455 -2390 -449
rect -2448 -489 -2436 -455
rect -2402 -489 -2390 -455
rect -2448 -495 -2390 -489
rect -2330 -455 -2272 -449
rect -2330 -489 -2318 -455
rect -2284 -489 -2272 -455
rect -2330 -495 -2272 -489
rect -2212 -455 -2154 -449
rect -2212 -489 -2200 -455
rect -2166 -489 -2154 -455
rect -2212 -495 -2154 -489
rect -2094 -455 -2036 -449
rect -2094 -489 -2082 -455
rect -2048 -489 -2036 -455
rect -2094 -495 -2036 -489
rect -1976 -455 -1918 -449
rect -1976 -489 -1964 -455
rect -1930 -489 -1918 -455
rect -1976 -495 -1918 -489
rect -1858 -455 -1800 -449
rect -1858 -489 -1846 -455
rect -1812 -489 -1800 -455
rect -1858 -495 -1800 -489
rect -1740 -455 -1682 -449
rect -1740 -489 -1728 -455
rect -1694 -489 -1682 -455
rect -1740 -495 -1682 -489
rect -1622 -455 -1564 -449
rect -1622 -489 -1610 -455
rect -1576 -489 -1564 -455
rect -1622 -495 -1564 -489
rect -1504 -455 -1446 -449
rect -1504 -489 -1492 -455
rect -1458 -489 -1446 -455
rect -1504 -495 -1446 -489
rect -1386 -455 -1328 -449
rect -1386 -489 -1374 -455
rect -1340 -489 -1328 -455
rect -1386 -495 -1328 -489
rect -1268 -455 -1210 -449
rect -1268 -489 -1256 -455
rect -1222 -489 -1210 -455
rect -1268 -495 -1210 -489
rect -1150 -455 -1092 -449
rect -1150 -489 -1138 -455
rect -1104 -489 -1092 -455
rect -1150 -495 -1092 -489
rect -1032 -455 -974 -449
rect -1032 -489 -1020 -455
rect -986 -489 -974 -455
rect -1032 -495 -974 -489
rect -914 -455 -856 -449
rect -914 -489 -902 -455
rect -868 -489 -856 -455
rect -914 -495 -856 -489
rect -796 -455 -738 -449
rect -796 -489 -784 -455
rect -750 -489 -738 -455
rect -796 -495 -738 -489
rect -678 -455 -620 -449
rect -678 -489 -666 -455
rect -632 -489 -620 -455
rect -678 -495 -620 -489
rect -560 -455 -502 -449
rect -560 -489 -548 -455
rect -514 -489 -502 -455
rect -560 -495 -502 -489
rect -442 -455 -384 -449
rect -442 -489 -430 -455
rect -396 -489 -384 -455
rect -442 -495 -384 -489
rect -324 -455 -266 -449
rect -324 -489 -312 -455
rect -278 -489 -266 -455
rect -324 -495 -266 -489
rect -206 -455 -148 -449
rect -206 -489 -194 -455
rect -160 -489 -148 -455
rect -206 -495 -148 -489
rect -88 -455 -30 -449
rect -88 -489 -76 -455
rect -42 -489 -30 -455
rect -88 -495 -30 -489
rect 30 -455 88 -449
rect 30 -489 42 -455
rect 76 -489 88 -455
rect 30 -495 88 -489
rect 148 -455 206 -449
rect 148 -489 160 -455
rect 194 -489 206 -455
rect 148 -495 206 -489
rect 266 -455 324 -449
rect 266 -489 278 -455
rect 312 -489 324 -455
rect 266 -495 324 -489
rect 384 -455 442 -449
rect 384 -489 396 -455
rect 430 -489 442 -455
rect 384 -495 442 -489
rect 502 -455 560 -449
rect 502 -489 514 -455
rect 548 -489 560 -455
rect 502 -495 560 -489
rect 620 -455 678 -449
rect 620 -489 632 -455
rect 666 -489 678 -455
rect 620 -495 678 -489
rect 738 -455 796 -449
rect 738 -489 750 -455
rect 784 -489 796 -455
rect 738 -495 796 -489
rect 856 -455 914 -449
rect 856 -489 868 -455
rect 902 -489 914 -455
rect 856 -495 914 -489
rect 974 -455 1032 -449
rect 974 -489 986 -455
rect 1020 -489 1032 -455
rect 974 -495 1032 -489
rect 1092 -455 1150 -449
rect 1092 -489 1104 -455
rect 1138 -489 1150 -455
rect 1092 -495 1150 -489
rect 1210 -455 1268 -449
rect 1210 -489 1222 -455
rect 1256 -489 1268 -455
rect 1210 -495 1268 -489
rect 1328 -455 1386 -449
rect 1328 -489 1340 -455
rect 1374 -489 1386 -455
rect 1328 -495 1386 -489
rect 1446 -455 1504 -449
rect 1446 -489 1458 -455
rect 1492 -489 1504 -455
rect 1446 -495 1504 -489
rect 1564 -455 1622 -449
rect 1564 -489 1576 -455
rect 1610 -489 1622 -455
rect 1564 -495 1622 -489
rect 1682 -455 1740 -449
rect 1682 -489 1694 -455
rect 1728 -489 1740 -455
rect 1682 -495 1740 -489
rect 1800 -455 1858 -449
rect 1800 -489 1812 -455
rect 1846 -489 1858 -455
rect 1800 -495 1858 -489
rect 1918 -455 1976 -449
rect 1918 -489 1930 -455
rect 1964 -489 1976 -455
rect 1918 -495 1976 -489
rect 2036 -455 2094 -449
rect 2036 -489 2048 -455
rect 2082 -489 2094 -455
rect 2036 -495 2094 -489
rect 2154 -455 2212 -449
rect 2154 -489 2166 -455
rect 2200 -489 2212 -455
rect 2154 -495 2212 -489
rect 2272 -455 2330 -449
rect 2272 -489 2284 -455
rect 2318 -489 2330 -455
rect 2272 -495 2330 -489
rect 2390 -455 2448 -449
rect 2390 -489 2402 -455
rect 2436 -489 2448 -455
rect 2390 -495 2448 -489
rect 2508 -455 2566 -449
rect 2508 -489 2520 -455
rect 2554 -489 2566 -455
rect 2508 -495 2566 -489
rect 2626 -455 2684 -449
rect 2626 -489 2638 -455
rect 2672 -489 2684 -455
rect 2626 -495 2684 -489
rect 2744 -455 2802 -449
rect 2744 -489 2756 -455
rect 2790 -489 2802 -455
rect 2744 -495 2802 -489
rect 2862 -455 2920 -449
rect 2862 -489 2874 -455
rect 2908 -489 2920 -455
rect 2862 -495 2920 -489
rect -2973 -548 -2927 -536
rect -2973 -1124 -2967 -548
rect -2933 -1124 -2927 -548
rect -2973 -1136 -2927 -1124
rect -2855 -548 -2809 -536
rect -2855 -1124 -2849 -548
rect -2815 -1124 -2809 -548
rect -2855 -1136 -2809 -1124
rect -2737 -548 -2691 -536
rect -2737 -1124 -2731 -548
rect -2697 -1124 -2691 -548
rect -2737 -1136 -2691 -1124
rect -2619 -548 -2573 -536
rect -2619 -1124 -2613 -548
rect -2579 -1124 -2573 -548
rect -2619 -1136 -2573 -1124
rect -2501 -548 -2455 -536
rect -2501 -1124 -2495 -548
rect -2461 -1124 -2455 -548
rect -2501 -1136 -2455 -1124
rect -2383 -548 -2337 -536
rect -2383 -1124 -2377 -548
rect -2343 -1124 -2337 -548
rect -2383 -1136 -2337 -1124
rect -2265 -548 -2219 -536
rect -2265 -1124 -2259 -548
rect -2225 -1124 -2219 -548
rect -2265 -1136 -2219 -1124
rect -2147 -548 -2101 -536
rect -2147 -1124 -2141 -548
rect -2107 -1124 -2101 -548
rect -2147 -1136 -2101 -1124
rect -2029 -548 -1983 -536
rect -2029 -1124 -2023 -548
rect -1989 -1124 -1983 -548
rect -2029 -1136 -1983 -1124
rect -1911 -548 -1865 -536
rect -1911 -1124 -1905 -548
rect -1871 -1124 -1865 -548
rect -1911 -1136 -1865 -1124
rect -1793 -548 -1747 -536
rect -1793 -1124 -1787 -548
rect -1753 -1124 -1747 -548
rect -1793 -1136 -1747 -1124
rect -1675 -548 -1629 -536
rect -1675 -1124 -1669 -548
rect -1635 -1124 -1629 -548
rect -1675 -1136 -1629 -1124
rect -1557 -548 -1511 -536
rect -1557 -1124 -1551 -548
rect -1517 -1124 -1511 -548
rect -1557 -1136 -1511 -1124
rect -1439 -548 -1393 -536
rect -1439 -1124 -1433 -548
rect -1399 -1124 -1393 -548
rect -1439 -1136 -1393 -1124
rect -1321 -548 -1275 -536
rect -1321 -1124 -1315 -548
rect -1281 -1124 -1275 -548
rect -1321 -1136 -1275 -1124
rect -1203 -548 -1157 -536
rect -1203 -1124 -1197 -548
rect -1163 -1124 -1157 -548
rect -1203 -1136 -1157 -1124
rect -1085 -548 -1039 -536
rect -1085 -1124 -1079 -548
rect -1045 -1124 -1039 -548
rect -1085 -1136 -1039 -1124
rect -967 -548 -921 -536
rect -967 -1124 -961 -548
rect -927 -1124 -921 -548
rect -967 -1136 -921 -1124
rect -849 -548 -803 -536
rect -849 -1124 -843 -548
rect -809 -1124 -803 -548
rect -849 -1136 -803 -1124
rect -731 -548 -685 -536
rect -731 -1124 -725 -548
rect -691 -1124 -685 -548
rect -731 -1136 -685 -1124
rect -613 -548 -567 -536
rect -613 -1124 -607 -548
rect -573 -1124 -567 -548
rect -613 -1136 -567 -1124
rect -495 -548 -449 -536
rect -495 -1124 -489 -548
rect -455 -1124 -449 -548
rect -495 -1136 -449 -1124
rect -377 -548 -331 -536
rect -377 -1124 -371 -548
rect -337 -1124 -331 -548
rect -377 -1136 -331 -1124
rect -259 -548 -213 -536
rect -259 -1124 -253 -548
rect -219 -1124 -213 -548
rect -259 -1136 -213 -1124
rect -141 -548 -95 -536
rect -141 -1124 -135 -548
rect -101 -1124 -95 -548
rect -141 -1136 -95 -1124
rect -23 -548 23 -536
rect -23 -1124 -17 -548
rect 17 -1124 23 -548
rect -23 -1136 23 -1124
rect 95 -548 141 -536
rect 95 -1124 101 -548
rect 135 -1124 141 -548
rect 95 -1136 141 -1124
rect 213 -548 259 -536
rect 213 -1124 219 -548
rect 253 -1124 259 -548
rect 213 -1136 259 -1124
rect 331 -548 377 -536
rect 331 -1124 337 -548
rect 371 -1124 377 -548
rect 331 -1136 377 -1124
rect 449 -548 495 -536
rect 449 -1124 455 -548
rect 489 -1124 495 -548
rect 449 -1136 495 -1124
rect 567 -548 613 -536
rect 567 -1124 573 -548
rect 607 -1124 613 -548
rect 567 -1136 613 -1124
rect 685 -548 731 -536
rect 685 -1124 691 -548
rect 725 -1124 731 -548
rect 685 -1136 731 -1124
rect 803 -548 849 -536
rect 803 -1124 809 -548
rect 843 -1124 849 -548
rect 803 -1136 849 -1124
rect 921 -548 967 -536
rect 921 -1124 927 -548
rect 961 -1124 967 -548
rect 921 -1136 967 -1124
rect 1039 -548 1085 -536
rect 1039 -1124 1045 -548
rect 1079 -1124 1085 -548
rect 1039 -1136 1085 -1124
rect 1157 -548 1203 -536
rect 1157 -1124 1163 -548
rect 1197 -1124 1203 -548
rect 1157 -1136 1203 -1124
rect 1275 -548 1321 -536
rect 1275 -1124 1281 -548
rect 1315 -1124 1321 -548
rect 1275 -1136 1321 -1124
rect 1393 -548 1439 -536
rect 1393 -1124 1399 -548
rect 1433 -1124 1439 -548
rect 1393 -1136 1439 -1124
rect 1511 -548 1557 -536
rect 1511 -1124 1517 -548
rect 1551 -1124 1557 -548
rect 1511 -1136 1557 -1124
rect 1629 -548 1675 -536
rect 1629 -1124 1635 -548
rect 1669 -1124 1675 -548
rect 1629 -1136 1675 -1124
rect 1747 -548 1793 -536
rect 1747 -1124 1753 -548
rect 1787 -1124 1793 -548
rect 1747 -1136 1793 -1124
rect 1865 -548 1911 -536
rect 1865 -1124 1871 -548
rect 1905 -1124 1911 -548
rect 1865 -1136 1911 -1124
rect 1983 -548 2029 -536
rect 1983 -1124 1989 -548
rect 2023 -1124 2029 -548
rect 1983 -1136 2029 -1124
rect 2101 -548 2147 -536
rect 2101 -1124 2107 -548
rect 2141 -1124 2147 -548
rect 2101 -1136 2147 -1124
rect 2219 -548 2265 -536
rect 2219 -1124 2225 -548
rect 2259 -1124 2265 -548
rect 2219 -1136 2265 -1124
rect 2337 -548 2383 -536
rect 2337 -1124 2343 -548
rect 2377 -1124 2383 -548
rect 2337 -1136 2383 -1124
rect 2455 -548 2501 -536
rect 2455 -1124 2461 -548
rect 2495 -1124 2501 -548
rect 2455 -1136 2501 -1124
rect 2573 -548 2619 -536
rect 2573 -1124 2579 -548
rect 2613 -1124 2619 -548
rect 2573 -1136 2619 -1124
rect 2691 -548 2737 -536
rect 2691 -1124 2697 -548
rect 2731 -1124 2737 -548
rect 2691 -1136 2737 -1124
rect 2809 -548 2855 -536
rect 2809 -1124 2815 -548
rect 2849 -1124 2855 -548
rect 2809 -1136 2855 -1124
rect 2927 -548 2973 -536
rect 2927 -1124 2933 -548
rect 2967 -1124 2973 -548
rect 2927 -1136 2973 -1124
rect -2920 -1183 -2862 -1177
rect -2920 -1217 -2908 -1183
rect -2874 -1217 -2862 -1183
rect -2920 -1223 -2862 -1217
rect -2802 -1183 -2744 -1177
rect -2802 -1217 -2790 -1183
rect -2756 -1217 -2744 -1183
rect -2802 -1223 -2744 -1217
rect -2684 -1183 -2626 -1177
rect -2684 -1217 -2672 -1183
rect -2638 -1217 -2626 -1183
rect -2684 -1223 -2626 -1217
rect -2566 -1183 -2508 -1177
rect -2566 -1217 -2554 -1183
rect -2520 -1217 -2508 -1183
rect -2566 -1223 -2508 -1217
rect -2448 -1183 -2390 -1177
rect -2448 -1217 -2436 -1183
rect -2402 -1217 -2390 -1183
rect -2448 -1223 -2390 -1217
rect -2330 -1183 -2272 -1177
rect -2330 -1217 -2318 -1183
rect -2284 -1217 -2272 -1183
rect -2330 -1223 -2272 -1217
rect -2212 -1183 -2154 -1177
rect -2212 -1217 -2200 -1183
rect -2166 -1217 -2154 -1183
rect -2212 -1223 -2154 -1217
rect -2094 -1183 -2036 -1177
rect -2094 -1217 -2082 -1183
rect -2048 -1217 -2036 -1183
rect -2094 -1223 -2036 -1217
rect -1976 -1183 -1918 -1177
rect -1976 -1217 -1964 -1183
rect -1930 -1217 -1918 -1183
rect -1976 -1223 -1918 -1217
rect -1858 -1183 -1800 -1177
rect -1858 -1217 -1846 -1183
rect -1812 -1217 -1800 -1183
rect -1858 -1223 -1800 -1217
rect -1740 -1183 -1682 -1177
rect -1740 -1217 -1728 -1183
rect -1694 -1217 -1682 -1183
rect -1740 -1223 -1682 -1217
rect -1622 -1183 -1564 -1177
rect -1622 -1217 -1610 -1183
rect -1576 -1217 -1564 -1183
rect -1622 -1223 -1564 -1217
rect -1504 -1183 -1446 -1177
rect -1504 -1217 -1492 -1183
rect -1458 -1217 -1446 -1183
rect -1504 -1223 -1446 -1217
rect -1386 -1183 -1328 -1177
rect -1386 -1217 -1374 -1183
rect -1340 -1217 -1328 -1183
rect -1386 -1223 -1328 -1217
rect -1268 -1183 -1210 -1177
rect -1268 -1217 -1256 -1183
rect -1222 -1217 -1210 -1183
rect -1268 -1223 -1210 -1217
rect -1150 -1183 -1092 -1177
rect -1150 -1217 -1138 -1183
rect -1104 -1217 -1092 -1183
rect -1150 -1223 -1092 -1217
rect -1032 -1183 -974 -1177
rect -1032 -1217 -1020 -1183
rect -986 -1217 -974 -1183
rect -1032 -1223 -974 -1217
rect -914 -1183 -856 -1177
rect -914 -1217 -902 -1183
rect -868 -1217 -856 -1183
rect -914 -1223 -856 -1217
rect -796 -1183 -738 -1177
rect -796 -1217 -784 -1183
rect -750 -1217 -738 -1183
rect -796 -1223 -738 -1217
rect -678 -1183 -620 -1177
rect -678 -1217 -666 -1183
rect -632 -1217 -620 -1183
rect -678 -1223 -620 -1217
rect -560 -1183 -502 -1177
rect -560 -1217 -548 -1183
rect -514 -1217 -502 -1183
rect -560 -1223 -502 -1217
rect -442 -1183 -384 -1177
rect -442 -1217 -430 -1183
rect -396 -1217 -384 -1183
rect -442 -1223 -384 -1217
rect -324 -1183 -266 -1177
rect -324 -1217 -312 -1183
rect -278 -1217 -266 -1183
rect -324 -1223 -266 -1217
rect -206 -1183 -148 -1177
rect -206 -1217 -194 -1183
rect -160 -1217 -148 -1183
rect -206 -1223 -148 -1217
rect -88 -1183 -30 -1177
rect -88 -1217 -76 -1183
rect -42 -1217 -30 -1183
rect -88 -1223 -30 -1217
rect 30 -1183 88 -1177
rect 30 -1217 42 -1183
rect 76 -1217 88 -1183
rect 30 -1223 88 -1217
rect 148 -1183 206 -1177
rect 148 -1217 160 -1183
rect 194 -1217 206 -1183
rect 148 -1223 206 -1217
rect 266 -1183 324 -1177
rect 266 -1217 278 -1183
rect 312 -1217 324 -1183
rect 266 -1223 324 -1217
rect 384 -1183 442 -1177
rect 384 -1217 396 -1183
rect 430 -1217 442 -1183
rect 384 -1223 442 -1217
rect 502 -1183 560 -1177
rect 502 -1217 514 -1183
rect 548 -1217 560 -1183
rect 502 -1223 560 -1217
rect 620 -1183 678 -1177
rect 620 -1217 632 -1183
rect 666 -1217 678 -1183
rect 620 -1223 678 -1217
rect 738 -1183 796 -1177
rect 738 -1217 750 -1183
rect 784 -1217 796 -1183
rect 738 -1223 796 -1217
rect 856 -1183 914 -1177
rect 856 -1217 868 -1183
rect 902 -1217 914 -1183
rect 856 -1223 914 -1217
rect 974 -1183 1032 -1177
rect 974 -1217 986 -1183
rect 1020 -1217 1032 -1183
rect 974 -1223 1032 -1217
rect 1092 -1183 1150 -1177
rect 1092 -1217 1104 -1183
rect 1138 -1217 1150 -1183
rect 1092 -1223 1150 -1217
rect 1210 -1183 1268 -1177
rect 1210 -1217 1222 -1183
rect 1256 -1217 1268 -1183
rect 1210 -1223 1268 -1217
rect 1328 -1183 1386 -1177
rect 1328 -1217 1340 -1183
rect 1374 -1217 1386 -1183
rect 1328 -1223 1386 -1217
rect 1446 -1183 1504 -1177
rect 1446 -1217 1458 -1183
rect 1492 -1217 1504 -1183
rect 1446 -1223 1504 -1217
rect 1564 -1183 1622 -1177
rect 1564 -1217 1576 -1183
rect 1610 -1217 1622 -1183
rect 1564 -1223 1622 -1217
rect 1682 -1183 1740 -1177
rect 1682 -1217 1694 -1183
rect 1728 -1217 1740 -1183
rect 1682 -1223 1740 -1217
rect 1800 -1183 1858 -1177
rect 1800 -1217 1812 -1183
rect 1846 -1217 1858 -1183
rect 1800 -1223 1858 -1217
rect 1918 -1183 1976 -1177
rect 1918 -1217 1930 -1183
rect 1964 -1217 1976 -1183
rect 1918 -1223 1976 -1217
rect 2036 -1183 2094 -1177
rect 2036 -1217 2048 -1183
rect 2082 -1217 2094 -1183
rect 2036 -1223 2094 -1217
rect 2154 -1183 2212 -1177
rect 2154 -1217 2166 -1183
rect 2200 -1217 2212 -1183
rect 2154 -1223 2212 -1217
rect 2272 -1183 2330 -1177
rect 2272 -1217 2284 -1183
rect 2318 -1217 2330 -1183
rect 2272 -1223 2330 -1217
rect 2390 -1183 2448 -1177
rect 2390 -1217 2402 -1183
rect 2436 -1217 2448 -1183
rect 2390 -1223 2448 -1217
rect 2508 -1183 2566 -1177
rect 2508 -1217 2520 -1183
rect 2554 -1217 2566 -1183
rect 2508 -1223 2566 -1217
rect 2626 -1183 2684 -1177
rect 2626 -1217 2638 -1183
rect 2672 -1217 2684 -1183
rect 2626 -1223 2684 -1217
rect 2744 -1183 2802 -1177
rect 2744 -1217 2756 -1183
rect 2790 -1217 2802 -1183
rect 2744 -1223 2802 -1217
rect 2862 -1183 2920 -1177
rect 2862 -1217 2874 -1183
rect 2908 -1217 2920 -1183
rect 2862 -1223 2920 -1217
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -3064 -1302 3064 1302
string parameters w 3 l 0.3 m 3 nf 50 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
