magic
tech sky130B
magscale 1 2
timestamp 1608096578
<< pwell >>
rect -701 -937 701 937
<< nmos >>
rect -505 527 -385 727
rect -327 527 -207 727
rect -149 527 -29 727
rect 29 527 149 727
rect 207 527 327 727
rect 385 527 505 727
rect -505 109 -385 309
rect -327 109 -207 309
rect -149 109 -29 309
rect 29 109 149 309
rect 207 109 327 309
rect 385 109 505 309
rect -505 -309 -385 -109
rect -327 -309 -207 -109
rect -149 -309 -29 -109
rect 29 -309 149 -109
rect 207 -309 327 -109
rect 385 -309 505 -109
rect -505 -727 -385 -527
rect -327 -727 -207 -527
rect -149 -727 -29 -527
rect 29 -727 149 -527
rect 207 -727 327 -527
rect 385 -727 505 -527
<< ndiff >>
rect -563 715 -505 727
rect -563 539 -551 715
rect -517 539 -505 715
rect -563 527 -505 539
rect -385 715 -327 727
rect -385 539 -373 715
rect -339 539 -327 715
rect -385 527 -327 539
rect -207 715 -149 727
rect -207 539 -195 715
rect -161 539 -149 715
rect -207 527 -149 539
rect -29 715 29 727
rect -29 539 -17 715
rect 17 539 29 715
rect -29 527 29 539
rect 149 715 207 727
rect 149 539 161 715
rect 195 539 207 715
rect 149 527 207 539
rect 327 715 385 727
rect 327 539 339 715
rect 373 539 385 715
rect 327 527 385 539
rect 505 715 563 727
rect 505 539 517 715
rect 551 539 563 715
rect 505 527 563 539
rect -563 297 -505 309
rect -563 121 -551 297
rect -517 121 -505 297
rect -563 109 -505 121
rect -385 297 -327 309
rect -385 121 -373 297
rect -339 121 -327 297
rect -385 109 -327 121
rect -207 297 -149 309
rect -207 121 -195 297
rect -161 121 -149 297
rect -207 109 -149 121
rect -29 297 29 309
rect -29 121 -17 297
rect 17 121 29 297
rect -29 109 29 121
rect 149 297 207 309
rect 149 121 161 297
rect 195 121 207 297
rect 149 109 207 121
rect 327 297 385 309
rect 327 121 339 297
rect 373 121 385 297
rect 327 109 385 121
rect 505 297 563 309
rect 505 121 517 297
rect 551 121 563 297
rect 505 109 563 121
rect -563 -121 -505 -109
rect -563 -297 -551 -121
rect -517 -297 -505 -121
rect -563 -309 -505 -297
rect -385 -121 -327 -109
rect -385 -297 -373 -121
rect -339 -297 -327 -121
rect -385 -309 -327 -297
rect -207 -121 -149 -109
rect -207 -297 -195 -121
rect -161 -297 -149 -121
rect -207 -309 -149 -297
rect -29 -121 29 -109
rect -29 -297 -17 -121
rect 17 -297 29 -121
rect -29 -309 29 -297
rect 149 -121 207 -109
rect 149 -297 161 -121
rect 195 -297 207 -121
rect 149 -309 207 -297
rect 327 -121 385 -109
rect 327 -297 339 -121
rect 373 -297 385 -121
rect 327 -309 385 -297
rect 505 -121 563 -109
rect 505 -297 517 -121
rect 551 -297 563 -121
rect 505 -309 563 -297
rect -563 -539 -505 -527
rect -563 -715 -551 -539
rect -517 -715 -505 -539
rect -563 -727 -505 -715
rect -385 -539 -327 -527
rect -385 -715 -373 -539
rect -339 -715 -327 -539
rect -385 -727 -327 -715
rect -207 -539 -149 -527
rect -207 -715 -195 -539
rect -161 -715 -149 -539
rect -207 -727 -149 -715
rect -29 -539 29 -527
rect -29 -715 -17 -539
rect 17 -715 29 -539
rect -29 -727 29 -715
rect 149 -539 207 -527
rect 149 -715 161 -539
rect 195 -715 207 -539
rect 149 -727 207 -715
rect 327 -539 385 -527
rect 327 -715 339 -539
rect 373 -715 385 -539
rect 327 -727 385 -715
rect 505 -539 563 -527
rect 505 -715 517 -539
rect 551 -715 563 -539
rect 505 -727 563 -715
<< ndiffc >>
rect -551 539 -517 715
rect -373 539 -339 715
rect -195 539 -161 715
rect -17 539 17 715
rect 161 539 195 715
rect 339 539 373 715
rect 517 539 551 715
rect -551 121 -517 297
rect -373 121 -339 297
rect -195 121 -161 297
rect -17 121 17 297
rect 161 121 195 297
rect 339 121 373 297
rect 517 121 551 297
rect -551 -297 -517 -121
rect -373 -297 -339 -121
rect -195 -297 -161 -121
rect -17 -297 17 -121
rect 161 -297 195 -121
rect 339 -297 373 -121
rect 517 -297 551 -121
rect -551 -715 -517 -539
rect -373 -715 -339 -539
rect -195 -715 -161 -539
rect -17 -715 17 -539
rect 161 -715 195 -539
rect 339 -715 373 -539
rect 517 -715 551 -539
<< psubdiff >>
rect -665 867 -569 901
rect 569 867 665 901
rect -665 805 -631 867
rect 631 805 665 867
rect -665 -867 -631 -805
rect 631 -867 665 -805
rect -665 -901 -569 -867
rect 569 -901 665 -867
<< psubdiffcont >>
rect -569 867 569 901
rect -665 -805 -631 805
rect 631 -805 665 805
rect -569 -901 569 -867
<< poly >>
rect -505 799 -385 815
rect -505 765 -489 799
rect -401 765 -385 799
rect -505 727 -385 765
rect -327 799 -207 815
rect -327 765 -311 799
rect -223 765 -207 799
rect -327 727 -207 765
rect -149 799 -29 815
rect -149 765 -133 799
rect -45 765 -29 799
rect -149 727 -29 765
rect 29 799 149 815
rect 29 765 45 799
rect 133 765 149 799
rect 29 727 149 765
rect 207 799 327 815
rect 207 765 223 799
rect 311 765 327 799
rect 207 727 327 765
rect 385 799 505 815
rect 385 765 401 799
rect 489 765 505 799
rect 385 727 505 765
rect -505 489 -385 527
rect -505 455 -489 489
rect -401 455 -385 489
rect -505 439 -385 455
rect -327 489 -207 527
rect -327 455 -311 489
rect -223 455 -207 489
rect -327 439 -207 455
rect -149 489 -29 527
rect -149 455 -133 489
rect -45 455 -29 489
rect -149 439 -29 455
rect 29 489 149 527
rect 29 455 45 489
rect 133 455 149 489
rect 29 439 149 455
rect 207 489 327 527
rect 207 455 223 489
rect 311 455 327 489
rect 207 439 327 455
rect 385 489 505 527
rect 385 455 401 489
rect 489 455 505 489
rect 385 439 505 455
rect -505 381 -385 397
rect -505 347 -489 381
rect -401 347 -385 381
rect -505 309 -385 347
rect -327 381 -207 397
rect -327 347 -311 381
rect -223 347 -207 381
rect -327 309 -207 347
rect -149 381 -29 397
rect -149 347 -133 381
rect -45 347 -29 381
rect -149 309 -29 347
rect 29 381 149 397
rect 29 347 45 381
rect 133 347 149 381
rect 29 309 149 347
rect 207 381 327 397
rect 207 347 223 381
rect 311 347 327 381
rect 207 309 327 347
rect 385 381 505 397
rect 385 347 401 381
rect 489 347 505 381
rect 385 309 505 347
rect -505 71 -385 109
rect -505 37 -489 71
rect -401 37 -385 71
rect -505 21 -385 37
rect -327 71 -207 109
rect -327 37 -311 71
rect -223 37 -207 71
rect -327 21 -207 37
rect -149 71 -29 109
rect -149 37 -133 71
rect -45 37 -29 71
rect -149 21 -29 37
rect 29 71 149 109
rect 29 37 45 71
rect 133 37 149 71
rect 29 21 149 37
rect 207 71 327 109
rect 207 37 223 71
rect 311 37 327 71
rect 207 21 327 37
rect 385 71 505 109
rect 385 37 401 71
rect 489 37 505 71
rect 385 21 505 37
rect -505 -37 -385 -21
rect -505 -71 -489 -37
rect -401 -71 -385 -37
rect -505 -109 -385 -71
rect -327 -37 -207 -21
rect -327 -71 -311 -37
rect -223 -71 -207 -37
rect -327 -109 -207 -71
rect -149 -37 -29 -21
rect -149 -71 -133 -37
rect -45 -71 -29 -37
rect -149 -109 -29 -71
rect 29 -37 149 -21
rect 29 -71 45 -37
rect 133 -71 149 -37
rect 29 -109 149 -71
rect 207 -37 327 -21
rect 207 -71 223 -37
rect 311 -71 327 -37
rect 207 -109 327 -71
rect 385 -37 505 -21
rect 385 -71 401 -37
rect 489 -71 505 -37
rect 385 -109 505 -71
rect -505 -347 -385 -309
rect -505 -381 -489 -347
rect -401 -381 -385 -347
rect -505 -397 -385 -381
rect -327 -347 -207 -309
rect -327 -381 -311 -347
rect -223 -381 -207 -347
rect -327 -397 -207 -381
rect -149 -347 -29 -309
rect -149 -381 -133 -347
rect -45 -381 -29 -347
rect -149 -397 -29 -381
rect 29 -347 149 -309
rect 29 -381 45 -347
rect 133 -381 149 -347
rect 29 -397 149 -381
rect 207 -347 327 -309
rect 207 -381 223 -347
rect 311 -381 327 -347
rect 207 -397 327 -381
rect 385 -347 505 -309
rect 385 -381 401 -347
rect 489 -381 505 -347
rect 385 -397 505 -381
rect -505 -455 -385 -439
rect -505 -489 -489 -455
rect -401 -489 -385 -455
rect -505 -527 -385 -489
rect -327 -455 -207 -439
rect -327 -489 -311 -455
rect -223 -489 -207 -455
rect -327 -527 -207 -489
rect -149 -455 -29 -439
rect -149 -489 -133 -455
rect -45 -489 -29 -455
rect -149 -527 -29 -489
rect 29 -455 149 -439
rect 29 -489 45 -455
rect 133 -489 149 -455
rect 29 -527 149 -489
rect 207 -455 327 -439
rect 207 -489 223 -455
rect 311 -489 327 -455
rect 207 -527 327 -489
rect 385 -455 505 -439
rect 385 -489 401 -455
rect 489 -489 505 -455
rect 385 -527 505 -489
rect -505 -765 -385 -727
rect -505 -799 -489 -765
rect -401 -799 -385 -765
rect -505 -815 -385 -799
rect -327 -765 -207 -727
rect -327 -799 -311 -765
rect -223 -799 -207 -765
rect -327 -815 -207 -799
rect -149 -765 -29 -727
rect -149 -799 -133 -765
rect -45 -799 -29 -765
rect -149 -815 -29 -799
rect 29 -765 149 -727
rect 29 -799 45 -765
rect 133 -799 149 -765
rect 29 -815 149 -799
rect 207 -765 327 -727
rect 207 -799 223 -765
rect 311 -799 327 -765
rect 207 -815 327 -799
rect 385 -765 505 -727
rect 385 -799 401 -765
rect 489 -799 505 -765
rect 385 -815 505 -799
<< polycont >>
rect -489 765 -401 799
rect -311 765 -223 799
rect -133 765 -45 799
rect 45 765 133 799
rect 223 765 311 799
rect 401 765 489 799
rect -489 455 -401 489
rect -311 455 -223 489
rect -133 455 -45 489
rect 45 455 133 489
rect 223 455 311 489
rect 401 455 489 489
rect -489 347 -401 381
rect -311 347 -223 381
rect -133 347 -45 381
rect 45 347 133 381
rect 223 347 311 381
rect 401 347 489 381
rect -489 37 -401 71
rect -311 37 -223 71
rect -133 37 -45 71
rect 45 37 133 71
rect 223 37 311 71
rect 401 37 489 71
rect -489 -71 -401 -37
rect -311 -71 -223 -37
rect -133 -71 -45 -37
rect 45 -71 133 -37
rect 223 -71 311 -37
rect 401 -71 489 -37
rect -489 -381 -401 -347
rect -311 -381 -223 -347
rect -133 -381 -45 -347
rect 45 -381 133 -347
rect 223 -381 311 -347
rect 401 -381 489 -347
rect -489 -489 -401 -455
rect -311 -489 -223 -455
rect -133 -489 -45 -455
rect 45 -489 133 -455
rect 223 -489 311 -455
rect 401 -489 489 -455
rect -489 -799 -401 -765
rect -311 -799 -223 -765
rect -133 -799 -45 -765
rect 45 -799 133 -765
rect 223 -799 311 -765
rect 401 -799 489 -765
<< locali >>
rect -665 867 -569 901
rect 569 867 665 901
rect -665 805 -631 867
rect 631 805 665 867
rect -505 765 -489 799
rect -401 765 -385 799
rect -327 765 -311 799
rect -223 765 -207 799
rect -149 765 -133 799
rect -45 765 -29 799
rect 29 765 45 799
rect 133 765 149 799
rect 207 765 223 799
rect 311 765 327 799
rect 385 765 401 799
rect 489 765 505 799
rect -551 715 -517 731
rect -551 523 -517 539
rect -373 715 -339 731
rect -373 523 -339 539
rect -195 715 -161 731
rect -195 523 -161 539
rect -17 715 17 731
rect -17 523 17 539
rect 161 715 195 731
rect 161 523 195 539
rect 339 715 373 731
rect 339 523 373 539
rect 517 715 551 731
rect 517 523 551 539
rect -505 455 -489 489
rect -401 455 -385 489
rect -327 455 -311 489
rect -223 455 -207 489
rect -149 455 -133 489
rect -45 455 -29 489
rect 29 455 45 489
rect 133 455 149 489
rect 207 455 223 489
rect 311 455 327 489
rect 385 455 401 489
rect 489 455 505 489
rect -505 347 -489 381
rect -401 347 -385 381
rect -327 347 -311 381
rect -223 347 -207 381
rect -149 347 -133 381
rect -45 347 -29 381
rect 29 347 45 381
rect 133 347 149 381
rect 207 347 223 381
rect 311 347 327 381
rect 385 347 401 381
rect 489 347 505 381
rect -551 297 -517 313
rect -551 105 -517 121
rect -373 297 -339 313
rect -373 105 -339 121
rect -195 297 -161 313
rect -195 105 -161 121
rect -17 297 17 313
rect -17 105 17 121
rect 161 297 195 313
rect 161 105 195 121
rect 339 297 373 313
rect 339 105 373 121
rect 517 297 551 313
rect 517 105 551 121
rect -505 37 -489 71
rect -401 37 -385 71
rect -327 37 -311 71
rect -223 37 -207 71
rect -149 37 -133 71
rect -45 37 -29 71
rect 29 37 45 71
rect 133 37 149 71
rect 207 37 223 71
rect 311 37 327 71
rect 385 37 401 71
rect 489 37 505 71
rect -505 -71 -489 -37
rect -401 -71 -385 -37
rect -327 -71 -311 -37
rect -223 -71 -207 -37
rect -149 -71 -133 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 133 -71 149 -37
rect 207 -71 223 -37
rect 311 -71 327 -37
rect 385 -71 401 -37
rect 489 -71 505 -37
rect -551 -121 -517 -105
rect -551 -313 -517 -297
rect -373 -121 -339 -105
rect -373 -313 -339 -297
rect -195 -121 -161 -105
rect -195 -313 -161 -297
rect -17 -121 17 -105
rect -17 -313 17 -297
rect 161 -121 195 -105
rect 161 -313 195 -297
rect 339 -121 373 -105
rect 339 -313 373 -297
rect 517 -121 551 -105
rect 517 -313 551 -297
rect -505 -381 -489 -347
rect -401 -381 -385 -347
rect -327 -381 -311 -347
rect -223 -381 -207 -347
rect -149 -381 -133 -347
rect -45 -381 -29 -347
rect 29 -381 45 -347
rect 133 -381 149 -347
rect 207 -381 223 -347
rect 311 -381 327 -347
rect 385 -381 401 -347
rect 489 -381 505 -347
rect -505 -489 -489 -455
rect -401 -489 -385 -455
rect -327 -489 -311 -455
rect -223 -489 -207 -455
rect -149 -489 -133 -455
rect -45 -489 -29 -455
rect 29 -489 45 -455
rect 133 -489 149 -455
rect 207 -489 223 -455
rect 311 -489 327 -455
rect 385 -489 401 -455
rect 489 -489 505 -455
rect -551 -539 -517 -523
rect -551 -731 -517 -715
rect -373 -539 -339 -523
rect -373 -731 -339 -715
rect -195 -539 -161 -523
rect -195 -731 -161 -715
rect -17 -539 17 -523
rect -17 -731 17 -715
rect 161 -539 195 -523
rect 161 -731 195 -715
rect 339 -539 373 -523
rect 339 -731 373 -715
rect 517 -539 551 -523
rect 517 -731 551 -715
rect -505 -799 -489 -765
rect -401 -799 -385 -765
rect -327 -799 -311 -765
rect -223 -799 -207 -765
rect -149 -799 -133 -765
rect -45 -799 -29 -765
rect 29 -799 45 -765
rect 133 -799 149 -765
rect 207 -799 223 -765
rect 311 -799 327 -765
rect 385 -799 401 -765
rect 489 -799 505 -765
rect -665 -867 -631 -805
rect 631 -867 665 -805
rect -665 -901 -569 -867
rect 569 -901 665 -867
<< viali >>
rect -489 765 -401 799
rect -311 765 -223 799
rect -133 765 -45 799
rect 45 765 133 799
rect 223 765 311 799
rect 401 765 489 799
rect -551 539 -517 715
rect -373 539 -339 715
rect -195 539 -161 715
rect -17 539 17 715
rect 161 539 195 715
rect 339 539 373 715
rect 517 539 551 715
rect -489 455 -401 489
rect -311 455 -223 489
rect -133 455 -45 489
rect 45 455 133 489
rect 223 455 311 489
rect 401 455 489 489
rect -489 347 -401 381
rect -311 347 -223 381
rect -133 347 -45 381
rect 45 347 133 381
rect 223 347 311 381
rect 401 347 489 381
rect -551 121 -517 297
rect -373 121 -339 297
rect -195 121 -161 297
rect -17 121 17 297
rect 161 121 195 297
rect 339 121 373 297
rect 517 121 551 297
rect -489 37 -401 71
rect -311 37 -223 71
rect -133 37 -45 71
rect 45 37 133 71
rect 223 37 311 71
rect 401 37 489 71
rect -489 -71 -401 -37
rect -311 -71 -223 -37
rect -133 -71 -45 -37
rect 45 -71 133 -37
rect 223 -71 311 -37
rect 401 -71 489 -37
rect -551 -297 -517 -121
rect -373 -297 -339 -121
rect -195 -297 -161 -121
rect -17 -297 17 -121
rect 161 -297 195 -121
rect 339 -297 373 -121
rect 517 -297 551 -121
rect -489 -381 -401 -347
rect -311 -381 -223 -347
rect -133 -381 -45 -347
rect 45 -381 133 -347
rect 223 -381 311 -347
rect 401 -381 489 -347
rect -489 -489 -401 -455
rect -311 -489 -223 -455
rect -133 -489 -45 -455
rect 45 -489 133 -455
rect 223 -489 311 -455
rect 401 -489 489 -455
rect -551 -715 -517 -539
rect -373 -715 -339 -539
rect -195 -715 -161 -539
rect -17 -715 17 -539
rect 161 -715 195 -539
rect 339 -715 373 -539
rect 517 -715 551 -539
rect -489 -799 -401 -765
rect -311 -799 -223 -765
rect -133 -799 -45 -765
rect 45 -799 133 -765
rect 223 -799 311 -765
rect 401 -799 489 -765
<< metal1 >>
rect -10253 17051 -10243 18231
rect -10188 17051 -10178 18231
rect -9899 17050 -9889 18230
rect -9834 17050 -9824 18230
rect -9540 17050 -9530 18230
rect -9475 17050 -9465 18230
rect -9186 17048 -9176 18228
rect -9121 17048 -9111 18228
rect -8830 17053 -8820 18233
rect -8765 17053 -8755 18233
rect -8474 17058 -8464 18238
rect -8409 17058 -8399 18238
rect -8117 17061 -8107 18241
rect -8052 17061 -8042 18241
rect -7764 17062 -7754 18242
rect -7699 17062 -7689 18242
rect -7404 17058 -7394 18238
rect -7339 17058 -7329 18238
rect -501 799 -389 805
rect -501 765 -489 799
rect -401 765 -389 799
rect -501 759 -389 765
rect -323 799 -211 805
rect -323 765 -311 799
rect -223 765 -211 799
rect -323 759 -211 765
rect -145 799 -33 805
rect -145 765 -133 799
rect -45 765 -33 799
rect -145 759 -33 765
rect 33 799 145 805
rect 33 765 45 799
rect 133 765 145 799
rect 33 759 145 765
rect 211 799 323 805
rect 211 765 223 799
rect 311 765 323 799
rect 211 759 323 765
rect 389 799 501 805
rect 389 765 401 799
rect 489 765 501 799
rect 389 759 501 765
rect -557 715 -511 727
rect -557 539 -551 715
rect -517 539 -511 715
rect -557 527 -511 539
rect -379 715 -333 727
rect -379 539 -373 715
rect -339 539 -333 715
rect -379 527 -333 539
rect -201 715 -155 727
rect -201 539 -195 715
rect -161 539 -155 715
rect -201 527 -155 539
rect -23 715 23 727
rect -23 539 -17 715
rect 17 539 23 715
rect -23 527 23 539
rect 155 715 201 727
rect 155 539 161 715
rect 195 539 201 715
rect 155 527 201 539
rect 333 715 379 727
rect 333 539 339 715
rect 373 539 379 715
rect 333 527 379 539
rect 511 715 557 727
rect 511 539 517 715
rect 551 539 557 715
rect 511 527 557 539
rect -501 489 -389 495
rect -501 455 -489 489
rect -401 455 -389 489
rect -501 449 -389 455
rect -323 489 -211 495
rect -323 455 -311 489
rect -223 455 -211 489
rect -323 449 -211 455
rect -145 489 -33 495
rect -145 455 -133 489
rect -45 455 -33 489
rect -145 449 -33 455
rect 33 489 145 495
rect 33 455 45 489
rect 133 455 145 489
rect 33 449 145 455
rect 211 489 323 495
rect 211 455 223 489
rect 311 455 323 489
rect 211 449 323 455
rect 389 489 501 495
rect 389 455 401 489
rect 489 455 501 489
rect 389 449 501 455
rect -501 381 -389 387
rect -501 347 -489 381
rect -401 347 -389 381
rect -501 341 -389 347
rect -323 381 -211 387
rect -323 347 -311 381
rect -223 347 -211 381
rect -323 341 -211 347
rect -145 381 -33 387
rect -145 347 -133 381
rect -45 347 -33 381
rect -145 341 -33 347
rect 33 381 145 387
rect 33 347 45 381
rect 133 347 145 381
rect 33 341 145 347
rect 211 381 323 387
rect 211 347 223 381
rect 311 347 323 381
rect 211 341 323 347
rect 389 381 501 387
rect 389 347 401 381
rect 489 347 501 381
rect 389 341 501 347
rect -557 297 -511 309
rect -557 121 -551 297
rect -517 121 -511 297
rect -557 109 -511 121
rect -379 297 -333 309
rect -379 121 -373 297
rect -339 121 -333 297
rect -379 109 -333 121
rect -201 297 -155 309
rect -201 121 -195 297
rect -161 121 -155 297
rect -201 109 -155 121
rect -23 297 23 309
rect -23 121 -17 297
rect 17 121 23 297
rect -23 109 23 121
rect 155 297 201 309
rect 155 121 161 297
rect 195 121 201 297
rect 155 109 201 121
rect 333 297 379 309
rect 333 121 339 297
rect 373 121 379 297
rect 333 109 379 121
rect 511 297 557 309
rect 511 121 517 297
rect 551 121 557 297
rect 511 109 557 121
rect -501 71 -389 77
rect -501 37 -489 71
rect -401 37 -389 71
rect -501 31 -389 37
rect -323 71 -211 77
rect -323 37 -311 71
rect -223 37 -211 71
rect -323 31 -211 37
rect -145 71 -33 77
rect -145 37 -133 71
rect -45 37 -33 71
rect -145 31 -33 37
rect 33 71 145 77
rect 33 37 45 71
rect 133 37 145 71
rect 33 31 145 37
rect 211 71 323 77
rect 211 37 223 71
rect 311 37 323 71
rect 211 31 323 37
rect 389 71 501 77
rect 389 37 401 71
rect 489 37 501 71
rect 389 31 501 37
rect -501 -37 -389 -31
rect -501 -71 -489 -37
rect -401 -71 -389 -37
rect -501 -77 -389 -71
rect -323 -37 -211 -31
rect -323 -71 -311 -37
rect -223 -71 -211 -37
rect -323 -77 -211 -71
rect -145 -37 -33 -31
rect -145 -71 -133 -37
rect -45 -71 -33 -37
rect -145 -77 -33 -71
rect 33 -37 145 -31
rect 33 -71 45 -37
rect 133 -71 145 -37
rect 33 -77 145 -71
rect 211 -37 323 -31
rect 211 -71 223 -37
rect 311 -71 323 -37
rect 211 -77 323 -71
rect 389 -37 501 -31
rect 389 -71 401 -37
rect 489 -71 501 -37
rect 389 -77 501 -71
rect -557 -121 -511 -109
rect -557 -297 -551 -121
rect -517 -297 -511 -121
rect -557 -309 -511 -297
rect -379 -121 -333 -109
rect -379 -297 -373 -121
rect -339 -297 -333 -121
rect -379 -309 -333 -297
rect -201 -121 -155 -109
rect -201 -297 -195 -121
rect -161 -297 -155 -121
rect -201 -309 -155 -297
rect -23 -121 23 -109
rect -23 -297 -17 -121
rect 17 -297 23 -121
rect -23 -309 23 -297
rect 155 -121 201 -109
rect 155 -297 161 -121
rect 195 -297 201 -121
rect 155 -309 201 -297
rect 333 -121 379 -109
rect 333 -297 339 -121
rect 373 -297 379 -121
rect 333 -309 379 -297
rect 511 -121 557 -109
rect 511 -297 517 -121
rect 551 -297 557 -121
rect 511 -309 557 -297
rect -501 -347 -389 -341
rect -501 -381 -489 -347
rect -401 -381 -389 -347
rect -501 -387 -389 -381
rect -323 -347 -211 -341
rect -323 -381 -311 -347
rect -223 -381 -211 -347
rect -323 -387 -211 -381
rect -145 -347 -33 -341
rect -145 -381 -133 -347
rect -45 -381 -33 -347
rect -145 -387 -33 -381
rect 33 -347 145 -341
rect 33 -381 45 -347
rect 133 -381 145 -347
rect 33 -387 145 -381
rect 211 -347 323 -341
rect 211 -381 223 -347
rect 311 -381 323 -347
rect 211 -387 323 -381
rect 389 -347 501 -341
rect 389 -381 401 -347
rect 489 -381 501 -347
rect 389 -387 501 -381
rect -501 -455 -389 -449
rect -501 -489 -489 -455
rect -401 -489 -389 -455
rect -501 -495 -389 -489
rect -323 -455 -211 -449
rect -323 -489 -311 -455
rect -223 -489 -211 -455
rect -323 -495 -211 -489
rect -145 -455 -33 -449
rect -145 -489 -133 -455
rect -45 -489 -33 -455
rect -145 -495 -33 -489
rect 33 -455 145 -449
rect 33 -489 45 -455
rect 133 -489 145 -455
rect 33 -495 145 -489
rect 211 -455 323 -449
rect 211 -489 223 -455
rect 311 -489 323 -455
rect 211 -495 323 -489
rect 389 -455 501 -449
rect 389 -489 401 -455
rect 489 -489 501 -455
rect 389 -495 501 -489
rect -557 -539 -511 -527
rect -557 -715 -551 -539
rect -517 -715 -511 -539
rect -557 -727 -511 -715
rect -379 -539 -333 -527
rect -379 -715 -373 -539
rect -339 -715 -333 -539
rect -379 -727 -333 -715
rect -201 -539 -155 -527
rect -201 -715 -195 -539
rect -161 -715 -155 -539
rect -201 -727 -155 -715
rect -23 -539 23 -527
rect -23 -715 -17 -539
rect 17 -715 23 -539
rect -23 -727 23 -715
rect 155 -539 201 -527
rect 155 -715 161 -539
rect 195 -715 201 -539
rect 155 -727 201 -715
rect 333 -539 379 -527
rect 333 -715 339 -539
rect 373 -715 379 -539
rect 333 -727 379 -715
rect 511 -539 557 -527
rect 511 -715 517 -539
rect 551 -715 557 -539
rect 511 -727 557 -715
rect -501 -765 -389 -759
rect -501 -799 -489 -765
rect -401 -799 -389 -765
rect -501 -805 -389 -799
rect -323 -765 -211 -759
rect -323 -799 -311 -765
rect -223 -799 -211 -765
rect -323 -805 -211 -799
rect -145 -765 -33 -759
rect -145 -799 -133 -765
rect -45 -799 -33 -765
rect -145 -805 -33 -799
rect 33 -765 145 -759
rect 33 -799 45 -765
rect 133 -799 145 -765
rect 33 -805 145 -799
rect 211 -765 323 -759
rect 211 -799 223 -765
rect 311 -799 323 -765
rect 211 -805 323 -799
rect 389 -765 501 -759
rect 389 -799 401 -765
rect 489 -799 501 -765
rect 389 -805 501 -799
<< via1 >>
rect -10243 17051 -10188 18231
rect -9889 17050 -9834 18230
rect -9530 17050 -9475 18230
rect -9176 17048 -9121 18228
rect -8820 17053 -8765 18233
rect -8464 17058 -8409 18238
rect -8107 17061 -8052 18241
rect -7754 17062 -7699 18242
rect -7394 17058 -7339 18238
<< metal2 >>
rect -10243 18231 -10188 18241
rect -10243 17041 -10188 17051
rect -9889 18230 -9834 18240
rect -9889 17040 -9834 17050
rect -9530 18230 -9475 18240
rect -9530 17040 -9475 17050
rect -9176 18228 -9121 18238
rect -9176 17038 -9121 17048
rect -8820 18233 -8765 18243
rect -8820 17043 -8765 17053
rect -8464 18238 -8409 18248
rect -8464 17048 -8409 17058
rect -8107 18241 -8052 18251
rect -8107 17051 -8052 17061
rect -7754 18242 -7699 18252
rect -7754 17052 -7699 17062
rect -7394 18238 -7339 18248
rect -7394 17048 -7339 17058
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -648 -884 648 884
string parameters w 1 l 0.6 m 4 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
