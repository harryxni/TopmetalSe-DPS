magic
tech sky130B
magscale 1 2
timestamp 1662163768
<< nwell >>
rect -275 3700 43445 4050
rect 2805 3640 3469 3700
<< metal1 >>
rect -300 170 6720 270
<< metal3 >>
rect -245 810 6855 880
rect -290 500 6820 560
use bottom_pixel  bottom_pixel_0
timestamp 1662163768
transform 1 0 470 0 1 7290
box -770 -7420 3480 640
use bottom_pixel  bottom_pixel_1
timestamp 1662163768
transform 1 0 3470 0 1 7290
box -770 -7420 3480 640
use bottom_pixel  bottom_pixel_2
timestamp 1662163768
transform 1 0 9470 0 1 7290
box -770 -7420 3480 640
use bottom_pixel  bottom_pixel_3
timestamp 1662163768
transform 1 0 6470 0 1 7290
box -770 -7420 3480 640
use bottom_pixel  bottom_pixel_4
timestamp 1662163768
transform 1 0 15470 0 1 7290
box -770 -7420 3480 640
use bottom_pixel  bottom_pixel_5
timestamp 1662163768
transform 1 0 12470 0 1 7290
box -770 -7420 3480 640
use bottom_pixel  bottom_pixel_6
timestamp 1662163768
transform 1 0 21470 0 1 7290
box -770 -7420 3480 640
use bottom_pixel  bottom_pixel_7
timestamp 1662163768
transform 1 0 18470 0 1 7290
box -770 -7420 3480 640
use bottom_pixel  bottom_pixel_8
timestamp 1662163768
transform 1 0 27470 0 1 7290
box -770 -7420 3480 640
use bottom_pixel  bottom_pixel_9
timestamp 1662163768
transform 1 0 24470 0 1 7290
box -770 -7420 3480 640
use bottom_pixel  bottom_pixel_10
timestamp 1662163768
transform 1 0 33470 0 1 7290
box -770 -7420 3480 640
use bottom_pixel  bottom_pixel_11
timestamp 1662163768
transform 1 0 30470 0 1 7290
box -770 -7420 3480 640
use bottom_pixel  bottom_pixel_12
timestamp 1662163768
transform 1 0 39470 0 1 7290
box -770 -7420 3480 640
use bottom_pixel  bottom_pixel_13
timestamp 1662163768
transform 1 0 36470 0 1 7290
box -770 -7420 3480 640
<< end >>
