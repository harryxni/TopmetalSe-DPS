magic
tech sky130B
magscale 1 2
timestamp 1607692587
<< nwell >>
rect 24 934 4132 1252
rect 24 872 1632 934
rect 392 846 1632 872
rect 460 816 1632 846
rect 482 806 1632 816
rect 2316 786 4132 934
rect 2316 778 3884 786
rect 2316 776 2576 778
rect 2316 716 2502 776
rect 120 234 630 336
rect 120 64 780 234
rect 2110 230 2278 320
rect 2110 62 2482 230
<< pwell >>
rect 288 662 374 702
rect 452 662 538 702
rect 616 662 702 702
rect 780 662 866 702
rect 942 662 1028 702
rect 1108 662 1194 702
rect 2444 572 2530 612
rect 2606 572 2692 612
rect 2774 572 2860 612
rect 2940 608 3026 612
rect 2938 574 3026 608
rect 2940 572 3026 574
rect 3100 572 3186 612
rect 3264 570 3350 610
rect 3418 572 3504 612
rect 3586 570 3672 610
rect 3748 572 3834 612
<< nmos >>
rect 1720 720 1804 750
rect 238 404 268 488
rect 486 404 516 488
rect 776 464 864 494
rect 924 464 1884 494
rect 2108 466 2192 496
rect 924 352 2004 382
<< pmos >>
rect 496 1130 4096 1160
rect 344 1032 432 1062
rect 496 1032 4096 1062
rect 496 920 1576 950
rect 2370 818 2454 848
rect 238 140 268 284
rect 486 140 516 284
rect 2146 188 2230 218
<< ndiff >>
rect 1720 800 1804 816
rect 1720 766 1746 800
rect 1780 766 1804 800
rect 1720 750 1804 766
rect 1720 704 1804 720
rect 1720 670 1746 704
rect 1780 670 1804 704
rect 1720 654 1804 670
rect 776 544 864 560
rect 776 510 802 544
rect 836 510 864 544
rect 776 494 864 510
rect 924 544 1884 560
rect 924 510 932 544
rect 966 510 1000 544
rect 1034 510 1068 544
rect 1102 510 1136 544
rect 1170 510 1204 544
rect 1238 510 1272 544
rect 1306 510 1340 544
rect 1374 510 1408 544
rect 1442 510 1476 544
rect 1510 510 1544 544
rect 1578 510 1612 544
rect 1646 510 1680 544
rect 1714 510 1748 544
rect 1782 510 1816 544
rect 1850 510 1884 544
rect 924 494 1884 510
rect 2108 546 2192 562
rect 2108 512 2140 546
rect 2174 512 2192 546
rect 2108 496 2192 512
rect 174 460 238 488
rect 174 426 188 460
rect 222 426 238 460
rect 174 404 238 426
rect 268 460 334 488
rect 268 426 284 460
rect 318 426 334 460
rect 268 404 334 426
rect 422 460 486 488
rect 422 426 436 460
rect 470 426 486 460
rect 422 404 486 426
rect 516 460 582 488
rect 516 426 532 460
rect 566 426 582 460
rect 516 404 582 426
rect 776 448 864 464
rect 776 414 802 448
rect 836 414 864 448
rect 776 398 864 414
rect 924 448 1884 464
rect 924 432 2004 448
rect 924 398 940 432
rect 974 398 1008 432
rect 1042 398 1076 432
rect 1110 398 1144 432
rect 1178 398 1212 432
rect 1246 398 1280 432
rect 1314 398 1348 432
rect 1382 398 1416 432
rect 1450 398 1484 432
rect 1518 398 1552 432
rect 1586 398 1620 432
rect 1654 398 1688 432
rect 1722 398 1756 432
rect 1790 398 1824 432
rect 1858 398 1892 432
rect 1926 398 2004 432
rect 2108 442 2192 466
rect 2108 408 2134 442
rect 2168 408 2192 442
rect 2108 400 2192 408
rect 924 382 2004 398
rect 924 336 2004 352
rect 924 302 940 336
rect 974 302 1008 336
rect 1042 302 1076 336
rect 1110 302 1144 336
rect 1178 302 1212 336
rect 1246 302 1280 336
rect 1314 302 1348 336
rect 1382 302 1416 336
rect 1450 302 1484 336
rect 1518 302 1552 336
rect 1586 302 1620 336
rect 1654 302 1688 336
rect 1722 302 1756 336
rect 1790 302 1824 336
rect 1858 302 1892 336
rect 1926 302 2004 336
rect 924 286 2004 302
<< pdiff >>
rect 496 1206 4096 1216
rect 496 1172 514 1206
rect 548 1172 582 1206
rect 616 1172 650 1206
rect 684 1172 718 1206
rect 752 1172 786 1206
rect 820 1172 854 1206
rect 888 1172 922 1206
rect 956 1172 990 1206
rect 1024 1172 1058 1206
rect 1092 1172 1126 1206
rect 1160 1172 1194 1206
rect 1228 1172 1262 1206
rect 1296 1172 1330 1206
rect 1364 1172 1398 1206
rect 1432 1172 1466 1206
rect 1500 1172 1534 1206
rect 1568 1172 1602 1206
rect 1636 1172 1670 1206
rect 1704 1172 1738 1206
rect 1772 1172 1806 1206
rect 1840 1172 1874 1206
rect 1908 1172 1942 1206
rect 1976 1172 2010 1206
rect 2044 1172 2078 1206
rect 2112 1172 2146 1206
rect 2180 1172 2214 1206
rect 2248 1172 2282 1206
rect 2316 1172 2350 1206
rect 2384 1172 2418 1206
rect 2452 1172 2486 1206
rect 2520 1172 2554 1206
rect 2588 1172 2622 1206
rect 2656 1172 2690 1206
rect 2724 1172 2758 1206
rect 2792 1172 2826 1206
rect 2860 1172 2894 1206
rect 2928 1172 2962 1206
rect 2996 1172 3030 1206
rect 3064 1172 3098 1206
rect 3132 1172 3166 1206
rect 3200 1172 3234 1206
rect 3268 1172 3302 1206
rect 3336 1172 3370 1206
rect 3404 1172 3438 1206
rect 3472 1172 3506 1206
rect 3540 1172 3574 1206
rect 3608 1172 3642 1206
rect 3676 1172 3710 1206
rect 3744 1172 3778 1206
rect 3812 1172 3846 1206
rect 3880 1172 3914 1206
rect 3948 1172 3982 1206
rect 4016 1172 4096 1206
rect 496 1160 4096 1172
rect 344 1114 432 1130
rect 344 1080 370 1114
rect 404 1080 432 1114
rect 344 1062 432 1080
rect 496 1114 4096 1130
rect 496 1080 514 1114
rect 548 1080 582 1114
rect 616 1080 650 1114
rect 684 1080 718 1114
rect 752 1080 786 1114
rect 820 1080 854 1114
rect 888 1080 922 1114
rect 956 1080 990 1114
rect 1024 1080 1058 1114
rect 1092 1080 1126 1114
rect 1160 1080 1194 1114
rect 1228 1080 1262 1114
rect 1296 1080 1330 1114
rect 1364 1080 1398 1114
rect 1432 1080 1466 1114
rect 1500 1080 1534 1114
rect 1568 1080 1602 1114
rect 1636 1080 1670 1114
rect 1704 1080 1738 1114
rect 1772 1080 1806 1114
rect 1840 1080 1874 1114
rect 1908 1080 1942 1114
rect 1976 1080 2010 1114
rect 2044 1080 2078 1114
rect 2112 1080 2146 1114
rect 2180 1080 2214 1114
rect 2248 1080 2282 1114
rect 2316 1080 2350 1114
rect 2384 1080 2418 1114
rect 2452 1080 2486 1114
rect 2520 1080 2554 1114
rect 2588 1080 2622 1114
rect 2656 1080 2690 1114
rect 2724 1080 2758 1114
rect 2792 1080 2826 1114
rect 2860 1080 2894 1114
rect 2928 1080 2962 1114
rect 2996 1080 3030 1114
rect 3064 1080 3098 1114
rect 3132 1080 3166 1114
rect 3200 1080 3234 1114
rect 3268 1080 3302 1114
rect 3336 1080 3370 1114
rect 3404 1080 3438 1114
rect 3472 1080 3506 1114
rect 3540 1080 3574 1114
rect 3608 1080 3642 1114
rect 3676 1080 3710 1114
rect 3744 1080 3778 1114
rect 3812 1080 3846 1114
rect 3880 1080 3914 1114
rect 3948 1080 3982 1114
rect 4016 1080 4096 1114
rect 496 1062 4096 1080
rect 344 1016 432 1032
rect 344 982 372 1016
rect 406 982 432 1016
rect 344 966 432 982
rect 496 1016 4096 1032
rect 496 982 514 1016
rect 548 982 582 1016
rect 616 982 650 1016
rect 684 982 718 1016
rect 752 982 786 1016
rect 820 982 854 1016
rect 888 982 922 1016
rect 956 982 990 1016
rect 1024 982 1058 1016
rect 1092 982 1126 1016
rect 1160 982 1194 1016
rect 1228 982 1262 1016
rect 1296 982 1330 1016
rect 1364 982 1398 1016
rect 1432 982 1466 1016
rect 1500 982 1534 1016
rect 1568 982 1602 1016
rect 1636 982 1670 1016
rect 1704 982 1738 1016
rect 1772 982 1806 1016
rect 1840 982 1874 1016
rect 1908 982 1942 1016
rect 1976 982 2010 1016
rect 2044 982 2078 1016
rect 2112 982 2146 1016
rect 2180 982 2214 1016
rect 2248 982 2282 1016
rect 2316 982 2350 1016
rect 2384 982 2418 1016
rect 2452 982 2486 1016
rect 2520 982 2554 1016
rect 2588 982 2622 1016
rect 2656 982 2690 1016
rect 2724 982 2758 1016
rect 2792 982 2826 1016
rect 2860 982 2894 1016
rect 2928 982 2962 1016
rect 2996 982 3030 1016
rect 3064 982 3098 1016
rect 3132 982 3166 1016
rect 3200 982 3234 1016
rect 3268 982 3302 1016
rect 3336 982 3370 1016
rect 3404 982 3438 1016
rect 3472 982 3506 1016
rect 3540 982 3574 1016
rect 3608 982 3642 1016
rect 3676 982 3710 1016
rect 3744 982 3778 1016
rect 3812 982 3846 1016
rect 3880 982 3914 1016
rect 3948 982 3982 1016
rect 4016 982 4096 1016
rect 496 970 4096 982
rect 496 950 1576 970
rect 496 904 1576 920
rect 496 870 514 904
rect 548 870 582 904
rect 616 870 650 904
rect 684 870 718 904
rect 752 870 786 904
rect 820 870 854 904
rect 888 870 922 904
rect 956 870 990 904
rect 1024 870 1058 904
rect 1092 870 1126 904
rect 1160 870 1194 904
rect 1228 870 1262 904
rect 1296 870 1330 904
rect 1364 870 1398 904
rect 1432 870 1466 904
rect 1500 870 1576 904
rect 496 854 1576 870
rect 2370 898 2454 914
rect 2370 864 2396 898
rect 2430 864 2454 898
rect 2370 848 2454 864
rect 2370 802 2454 818
rect 2370 768 2388 802
rect 2422 768 2454 802
rect 2370 752 2454 768
rect 172 254 238 284
rect 172 220 188 254
rect 222 220 238 254
rect 172 182 238 220
rect 172 148 188 182
rect 222 148 238 182
rect 172 140 238 148
rect 268 276 334 284
rect 268 242 284 276
rect 318 242 334 276
rect 268 208 334 242
rect 268 174 284 208
rect 318 174 334 208
rect 268 140 334 174
rect 420 256 486 284
rect 420 222 436 256
rect 470 222 486 256
rect 420 182 486 222
rect 420 148 436 182
rect 470 148 486 182
rect 420 140 486 148
rect 516 276 582 284
rect 516 242 532 276
rect 566 242 582 276
rect 516 208 582 242
rect 2146 268 2230 284
rect 516 174 532 208
rect 566 174 582 208
rect 516 140 582 174
rect 2146 234 2172 268
rect 2206 234 2230 268
rect 2146 218 2230 234
rect 2146 172 2230 188
rect 2146 138 2172 172
rect 2206 138 2230 172
rect 2146 122 2230 138
<< ndiffc >>
rect 1746 766 1780 800
rect 1746 670 1780 704
rect 802 510 836 544
rect 932 510 966 544
rect 1000 510 1034 544
rect 1068 510 1102 544
rect 1136 510 1170 544
rect 1204 510 1238 544
rect 1272 510 1306 544
rect 1340 510 1374 544
rect 1408 510 1442 544
rect 1476 510 1510 544
rect 1544 510 1578 544
rect 1612 510 1646 544
rect 1680 510 1714 544
rect 1748 510 1782 544
rect 1816 510 1850 544
rect 2140 512 2174 546
rect 188 426 222 460
rect 284 426 318 460
rect 436 426 470 460
rect 532 426 566 460
rect 802 414 836 448
rect 940 398 974 432
rect 1008 398 1042 432
rect 1076 398 1110 432
rect 1144 398 1178 432
rect 1212 398 1246 432
rect 1280 398 1314 432
rect 1348 398 1382 432
rect 1416 398 1450 432
rect 1484 398 1518 432
rect 1552 398 1586 432
rect 1620 398 1654 432
rect 1688 398 1722 432
rect 1756 398 1790 432
rect 1824 398 1858 432
rect 1892 398 1926 432
rect 2134 408 2168 442
rect 940 302 974 336
rect 1008 302 1042 336
rect 1076 302 1110 336
rect 1144 302 1178 336
rect 1212 302 1246 336
rect 1280 302 1314 336
rect 1348 302 1382 336
rect 1416 302 1450 336
rect 1484 302 1518 336
rect 1552 302 1586 336
rect 1620 302 1654 336
rect 1688 302 1722 336
rect 1756 302 1790 336
rect 1824 302 1858 336
rect 1892 302 1926 336
<< pdiffc >>
rect 514 1172 548 1206
rect 582 1172 616 1206
rect 650 1172 684 1206
rect 718 1172 752 1206
rect 786 1172 820 1206
rect 854 1172 888 1206
rect 922 1172 956 1206
rect 990 1172 1024 1206
rect 1058 1172 1092 1206
rect 1126 1172 1160 1206
rect 1194 1172 1228 1206
rect 1262 1172 1296 1206
rect 1330 1172 1364 1206
rect 1398 1172 1432 1206
rect 1466 1172 1500 1206
rect 1534 1172 1568 1206
rect 1602 1172 1636 1206
rect 1670 1172 1704 1206
rect 1738 1172 1772 1206
rect 1806 1172 1840 1206
rect 1874 1172 1908 1206
rect 1942 1172 1976 1206
rect 2010 1172 2044 1206
rect 2078 1172 2112 1206
rect 2146 1172 2180 1206
rect 2214 1172 2248 1206
rect 2282 1172 2316 1206
rect 2350 1172 2384 1206
rect 2418 1172 2452 1206
rect 2486 1172 2520 1206
rect 2554 1172 2588 1206
rect 2622 1172 2656 1206
rect 2690 1172 2724 1206
rect 2758 1172 2792 1206
rect 2826 1172 2860 1206
rect 2894 1172 2928 1206
rect 2962 1172 2996 1206
rect 3030 1172 3064 1206
rect 3098 1172 3132 1206
rect 3166 1172 3200 1206
rect 3234 1172 3268 1206
rect 3302 1172 3336 1206
rect 3370 1172 3404 1206
rect 3438 1172 3472 1206
rect 3506 1172 3540 1206
rect 3574 1172 3608 1206
rect 3642 1172 3676 1206
rect 3710 1172 3744 1206
rect 3778 1172 3812 1206
rect 3846 1172 3880 1206
rect 3914 1172 3948 1206
rect 3982 1172 4016 1206
rect 370 1080 404 1114
rect 514 1080 548 1114
rect 582 1080 616 1114
rect 650 1080 684 1114
rect 718 1080 752 1114
rect 786 1080 820 1114
rect 854 1080 888 1114
rect 922 1080 956 1114
rect 990 1080 1024 1114
rect 1058 1080 1092 1114
rect 1126 1080 1160 1114
rect 1194 1080 1228 1114
rect 1262 1080 1296 1114
rect 1330 1080 1364 1114
rect 1398 1080 1432 1114
rect 1466 1080 1500 1114
rect 1534 1080 1568 1114
rect 1602 1080 1636 1114
rect 1670 1080 1704 1114
rect 1738 1080 1772 1114
rect 1806 1080 1840 1114
rect 1874 1080 1908 1114
rect 1942 1080 1976 1114
rect 2010 1080 2044 1114
rect 2078 1080 2112 1114
rect 2146 1080 2180 1114
rect 2214 1080 2248 1114
rect 2282 1080 2316 1114
rect 2350 1080 2384 1114
rect 2418 1080 2452 1114
rect 2486 1080 2520 1114
rect 2554 1080 2588 1114
rect 2622 1080 2656 1114
rect 2690 1080 2724 1114
rect 2758 1080 2792 1114
rect 2826 1080 2860 1114
rect 2894 1080 2928 1114
rect 2962 1080 2996 1114
rect 3030 1080 3064 1114
rect 3098 1080 3132 1114
rect 3166 1080 3200 1114
rect 3234 1080 3268 1114
rect 3302 1080 3336 1114
rect 3370 1080 3404 1114
rect 3438 1080 3472 1114
rect 3506 1080 3540 1114
rect 3574 1080 3608 1114
rect 3642 1080 3676 1114
rect 3710 1080 3744 1114
rect 3778 1080 3812 1114
rect 3846 1080 3880 1114
rect 3914 1080 3948 1114
rect 3982 1080 4016 1114
rect 372 982 406 1016
rect 514 982 548 1016
rect 582 982 616 1016
rect 650 982 684 1016
rect 718 982 752 1016
rect 786 982 820 1016
rect 854 982 888 1016
rect 922 982 956 1016
rect 990 982 1024 1016
rect 1058 982 1092 1016
rect 1126 982 1160 1016
rect 1194 982 1228 1016
rect 1262 982 1296 1016
rect 1330 982 1364 1016
rect 1398 982 1432 1016
rect 1466 982 1500 1016
rect 1534 982 1568 1016
rect 1602 982 1636 1016
rect 1670 982 1704 1016
rect 1738 982 1772 1016
rect 1806 982 1840 1016
rect 1874 982 1908 1016
rect 1942 982 1976 1016
rect 2010 982 2044 1016
rect 2078 982 2112 1016
rect 2146 982 2180 1016
rect 2214 982 2248 1016
rect 2282 982 2316 1016
rect 2350 982 2384 1016
rect 2418 982 2452 1016
rect 2486 982 2520 1016
rect 2554 982 2588 1016
rect 2622 982 2656 1016
rect 2690 982 2724 1016
rect 2758 982 2792 1016
rect 2826 982 2860 1016
rect 2894 982 2928 1016
rect 2962 982 2996 1016
rect 3030 982 3064 1016
rect 3098 982 3132 1016
rect 3166 982 3200 1016
rect 3234 982 3268 1016
rect 3302 982 3336 1016
rect 3370 982 3404 1016
rect 3438 982 3472 1016
rect 3506 982 3540 1016
rect 3574 982 3608 1016
rect 3642 982 3676 1016
rect 3710 982 3744 1016
rect 3778 982 3812 1016
rect 3846 982 3880 1016
rect 3914 982 3948 1016
rect 3982 982 4016 1016
rect 514 870 548 904
rect 582 870 616 904
rect 650 870 684 904
rect 718 870 752 904
rect 786 870 820 904
rect 854 870 888 904
rect 922 870 956 904
rect 990 870 1024 904
rect 1058 870 1092 904
rect 1126 870 1160 904
rect 1194 870 1228 904
rect 1262 870 1296 904
rect 1330 870 1364 904
rect 1398 870 1432 904
rect 1466 870 1500 904
rect 2396 864 2430 898
rect 2388 768 2422 802
rect 188 220 222 254
rect 188 148 222 182
rect 284 242 318 276
rect 284 174 318 208
rect 436 222 470 256
rect 436 148 470 182
rect 532 242 566 276
rect 532 174 566 208
rect 2172 234 2206 268
rect 2172 138 2206 172
<< psubdiff >>
rect 288 698 374 702
rect 288 664 314 698
rect 348 664 374 698
rect 288 662 374 664
rect 452 698 538 702
rect 452 664 478 698
rect 512 664 538 698
rect 452 662 538 664
rect 616 698 702 702
rect 616 664 642 698
rect 676 664 702 698
rect 616 662 702 664
rect 780 698 866 702
rect 780 664 806 698
rect 840 664 866 698
rect 780 662 866 664
rect 942 698 1028 702
rect 942 664 970 698
rect 1004 664 1028 698
rect 942 662 1028 664
rect 1108 698 1194 702
rect 1108 664 1134 698
rect 1168 664 1194 698
rect 1108 662 1194 664
rect 2444 608 2530 612
rect 2444 574 2470 608
rect 2504 574 2530 608
rect 2444 572 2530 574
rect 2606 608 2692 612
rect 2606 574 2634 608
rect 2668 574 2692 608
rect 2606 572 2692 574
rect 2774 608 2860 612
rect 2940 608 3026 612
rect 2774 574 2798 608
rect 2832 574 2860 608
rect 2938 574 2962 608
rect 2996 574 3026 608
rect 2774 572 2860 574
rect 2940 572 3026 574
rect 3100 608 3186 612
rect 3100 574 3126 608
rect 3160 574 3186 608
rect 3100 572 3186 574
rect 3264 608 3350 610
rect 3264 574 3290 608
rect 3324 574 3350 608
rect 3264 570 3350 574
rect 3418 608 3504 612
rect 3418 574 3446 608
rect 3480 574 3504 608
rect 3418 572 3504 574
rect 3586 608 3672 610
rect 3586 574 3610 608
rect 3644 574 3672 608
rect 3586 570 3672 574
rect 3748 608 3834 612
rect 3748 574 3774 608
rect 3808 574 3834 608
rect 3748 572 3834 574
<< nsubdiff >>
rect 2678 878 2760 880
rect 2678 844 2702 878
rect 2736 844 2760 878
rect 2678 842 2760 844
rect 2842 878 2924 880
rect 2842 844 2866 878
rect 2900 844 2924 878
rect 2842 842 2924 844
rect 3006 878 3088 880
rect 3006 844 3030 878
rect 3064 844 3088 878
rect 3006 842 3088 844
rect 3170 878 3252 880
rect 3170 844 3194 878
rect 3228 844 3252 878
rect 3170 842 3252 844
rect 3334 878 3416 880
rect 3334 844 3358 878
rect 3392 844 3416 878
rect 3334 842 3416 844
rect 3498 878 3580 880
rect 3498 844 3522 878
rect 3556 844 3580 878
rect 3498 842 3580 844
rect 3662 878 3744 880
rect 3662 844 3686 878
rect 3720 844 3744 878
rect 3662 842 3744 844
rect 3826 878 3908 880
rect 3826 844 3850 878
rect 3884 844 3908 878
rect 3826 842 3908 844
rect 662 134 744 138
rect 662 100 686 134
rect 720 100 744 134
rect 2336 156 2418 158
rect 2336 122 2360 156
rect 2394 122 2418 156
rect 2336 120 2418 122
<< psubdiffcont >>
rect 314 664 348 698
rect 478 664 512 698
rect 642 664 676 698
rect 806 664 840 698
rect 970 664 1004 698
rect 1134 664 1168 698
rect 2470 574 2504 608
rect 2634 574 2668 608
rect 2798 574 2832 608
rect 2962 574 2996 608
rect 3126 574 3160 608
rect 3290 574 3324 608
rect 3446 574 3480 608
rect 3610 574 3644 608
rect 3774 574 3808 608
<< nsubdiffcont >>
rect 2702 844 2736 878
rect 2866 844 2900 878
rect 3030 844 3064 878
rect 3194 844 3228 878
rect 3358 844 3392 878
rect 3522 844 3556 878
rect 3686 844 3720 878
rect 3850 844 3884 878
rect 686 100 720 134
rect 2360 122 2394 156
<< poly >>
rect 108 1160 480 1196
rect 108 1018 146 1160
rect 450 1130 496 1160
rect 4096 1130 4122 1160
rect 274 1032 344 1062
rect 432 1032 496 1062
rect 4096 1032 4122 1062
rect 260 1026 304 1032
rect 108 1002 196 1018
rect 108 968 138 1002
rect 172 968 196 1002
rect 250 1016 304 1026
rect 250 982 260 1016
rect 294 982 304 1016
rect 250 972 304 982
rect 108 954 196 968
rect 260 966 304 972
rect 438 920 496 950
rect 1576 920 1602 950
rect 438 866 472 920
rect 392 856 472 866
rect 392 822 408 856
rect 442 822 472 856
rect 392 812 472 822
rect 2244 850 2342 860
rect 2244 816 2260 850
rect 2294 848 2342 850
rect 2294 818 2370 848
rect 2454 818 2480 848
rect 2294 816 2342 818
rect 2244 806 2342 816
rect 1596 752 1650 768
rect 1596 718 1606 752
rect 1640 750 1650 752
rect 1640 720 1720 750
rect 1804 720 1830 750
rect 1640 718 1650 720
rect 1596 702 1650 718
rect 238 488 268 514
rect 486 488 516 514
rect 2004 548 2070 560
rect 2004 514 2020 548
rect 2054 514 2070 548
rect 2004 504 2070 514
rect 2034 496 2070 504
rect 704 464 776 494
rect 864 464 924 494
rect 1884 464 1914 494
rect 2034 466 2108 496
rect 2192 466 2218 496
rect 690 458 734 464
rect 680 448 734 458
rect 680 414 690 448
rect 724 414 734 448
rect 680 404 734 414
rect 238 376 268 404
rect 486 376 516 404
rect 690 398 734 404
rect 140 366 268 376
rect 140 332 156 366
rect 190 332 268 366
rect 140 322 268 332
rect 388 366 516 376
rect 388 332 404 366
rect 438 332 516 366
rect 850 352 924 382
rect 2004 352 2030 382
rect 850 342 898 352
rect 388 322 516 332
rect 238 284 268 322
rect 486 284 516 322
rect 800 329 898 342
rect 800 295 820 329
rect 854 295 898 329
rect 800 282 898 295
rect 2032 220 2086 236
rect 2032 186 2042 220
rect 2076 218 2086 220
rect 2076 188 2146 218
rect 2230 188 2256 218
rect 2076 186 2086 188
rect 2032 170 2086 186
rect 238 114 268 140
rect 486 114 516 140
<< polycont >>
rect 138 968 172 1002
rect 260 982 294 1016
rect 408 822 442 856
rect 2260 816 2294 850
rect 1606 718 1640 752
rect 2020 514 2054 548
rect 690 414 724 448
rect 156 332 190 366
rect 404 332 438 366
rect 820 295 854 329
rect 2042 186 2076 220
<< locali >>
rect 0 1214 42 1248
rect 76 1214 178 1248
rect 212 1214 314 1248
rect 348 1214 450 1248
rect 484 1214 586 1248
rect 620 1214 722 1248
rect 756 1214 858 1248
rect 892 1214 994 1248
rect 1028 1214 1130 1248
rect 1164 1214 1266 1248
rect 1300 1214 1402 1248
rect 1436 1214 1538 1248
rect 1572 1214 1674 1248
rect 1708 1214 1810 1248
rect 1844 1214 1946 1248
rect 1980 1214 2082 1248
rect 2116 1214 2218 1248
rect 2252 1214 2354 1248
rect 2388 1214 2490 1248
rect 2524 1214 2626 1248
rect 2660 1214 2762 1248
rect 2796 1214 2898 1248
rect 2932 1214 3034 1248
rect 3068 1214 3170 1248
rect 3204 1214 3306 1248
rect 3340 1214 3442 1248
rect 3476 1214 3578 1248
rect 3612 1214 3714 1248
rect 3748 1214 3850 1248
rect 3884 1214 3986 1248
rect 4020 1214 4132 1248
rect 496 1206 4096 1214
rect 496 1172 514 1206
rect 548 1172 582 1206
rect 616 1172 650 1206
rect 684 1172 718 1206
rect 752 1172 786 1206
rect 820 1172 854 1206
rect 888 1172 922 1206
rect 956 1172 990 1206
rect 1024 1172 1058 1206
rect 1092 1172 1126 1206
rect 1160 1172 1194 1206
rect 1228 1172 1262 1206
rect 1296 1172 1330 1206
rect 1364 1172 1398 1206
rect 1432 1172 1466 1206
rect 1500 1172 1534 1206
rect 1568 1172 1602 1206
rect 1636 1172 1670 1206
rect 1704 1172 1738 1206
rect 1772 1172 1806 1206
rect 1840 1172 1874 1206
rect 1908 1172 1942 1206
rect 1976 1172 2010 1206
rect 2044 1172 2078 1206
rect 2112 1172 2146 1206
rect 2180 1172 2214 1206
rect 2248 1172 2282 1206
rect 2316 1172 2350 1206
rect 2384 1172 2418 1206
rect 2452 1172 2486 1206
rect 2520 1172 2554 1206
rect 2588 1172 2622 1206
rect 2656 1172 2690 1206
rect 2724 1172 2758 1206
rect 2792 1172 2826 1206
rect 2860 1172 2894 1206
rect 2928 1172 2962 1206
rect 2996 1172 3030 1206
rect 3064 1172 3098 1206
rect 3132 1172 3166 1206
rect 3200 1172 3234 1206
rect 3268 1172 3302 1206
rect 3336 1172 3370 1206
rect 3404 1172 3438 1206
rect 3472 1172 3506 1206
rect 3540 1172 3574 1206
rect 3608 1172 3642 1206
rect 3676 1172 3710 1206
rect 3744 1172 3778 1206
rect 3812 1172 3846 1206
rect 3880 1172 3914 1206
rect 3948 1172 3982 1206
rect 4016 1172 4096 1206
rect 496 1170 4096 1172
rect 344 1114 4096 1116
rect 344 1080 370 1114
rect 404 1080 514 1114
rect 548 1080 582 1114
rect 616 1080 650 1114
rect 684 1080 718 1114
rect 752 1080 786 1114
rect 820 1080 854 1114
rect 888 1080 922 1114
rect 956 1080 990 1114
rect 1024 1080 1058 1114
rect 1092 1080 1126 1114
rect 1160 1080 1194 1114
rect 1228 1080 1262 1114
rect 1296 1080 1330 1114
rect 1364 1080 1398 1114
rect 1432 1080 1466 1114
rect 1500 1080 1534 1114
rect 1568 1080 1602 1114
rect 1636 1080 1670 1114
rect 1704 1080 1738 1114
rect 1772 1080 1806 1114
rect 1840 1080 1874 1114
rect 1908 1080 1942 1114
rect 1976 1080 2010 1114
rect 2044 1080 2078 1114
rect 2112 1080 2146 1114
rect 2180 1080 2214 1114
rect 2248 1080 2282 1114
rect 2316 1080 2350 1114
rect 2384 1080 2418 1114
rect 2452 1080 2486 1114
rect 2520 1080 2554 1114
rect 2596 1080 2622 1114
rect 2680 1080 2690 1114
rect 2724 1080 2758 1114
rect 2792 1080 2826 1114
rect 2860 1080 2894 1114
rect 2928 1080 2962 1114
rect 2996 1080 3030 1114
rect 3064 1080 3098 1114
rect 3132 1080 3166 1114
rect 3200 1080 3234 1114
rect 3268 1080 3302 1114
rect 3336 1080 3370 1114
rect 3404 1080 3438 1114
rect 3472 1080 3506 1114
rect 3540 1080 3574 1114
rect 3608 1080 3642 1114
rect 3676 1080 3710 1114
rect 3744 1080 3778 1114
rect 3812 1080 3846 1114
rect 3880 1080 3914 1114
rect 3948 1080 3982 1114
rect 4016 1080 4096 1114
rect 344 1078 4096 1080
rect 1674 1068 1750 1078
rect 1926 1068 2002 1078
rect 2374 1068 2450 1078
rect 244 1016 432 1018
rect 102 1002 192 1010
rect 102 968 138 1002
rect 172 968 192 1002
rect 244 982 260 1016
rect 294 982 372 1016
rect 406 982 432 1016
rect 244 980 432 982
rect 496 1016 4096 1018
rect 496 982 514 1016
rect 548 982 582 1016
rect 616 982 650 1016
rect 684 982 718 1016
rect 752 982 786 1016
rect 820 982 854 1016
rect 888 982 922 1016
rect 956 982 990 1016
rect 1024 982 1058 1016
rect 1092 982 1126 1016
rect 1160 982 1194 1016
rect 1228 982 1262 1016
rect 1296 982 1330 1016
rect 1364 982 1398 1016
rect 1432 982 1466 1016
rect 1500 982 1534 1016
rect 1568 982 1602 1016
rect 1636 982 1670 1016
rect 1704 982 1738 1016
rect 1772 982 1806 1016
rect 1840 982 1874 1016
rect 1908 982 1942 1016
rect 1976 982 2010 1016
rect 2044 982 2078 1016
rect 2112 982 2146 1016
rect 2180 982 2214 1016
rect 2248 982 2282 1016
rect 2316 982 2350 1016
rect 2384 982 2418 1016
rect 2452 982 2486 1016
rect 2520 982 2554 1016
rect 2588 982 2622 1016
rect 2656 982 2690 1016
rect 2724 982 2758 1016
rect 2792 982 2826 1016
rect 2860 982 2894 1016
rect 2928 982 2962 1016
rect 2996 982 3030 1016
rect 3064 982 3098 1016
rect 3132 982 3166 1016
rect 3200 982 3234 1016
rect 3268 982 3302 1016
rect 3336 982 3370 1016
rect 3404 982 3438 1016
rect 3472 982 3506 1016
rect 3540 982 3574 1016
rect 3608 982 3642 1016
rect 3676 982 3710 1016
rect 3744 982 3778 1016
rect 3812 982 3846 1016
rect 3880 982 3914 1016
rect 3948 982 3982 1016
rect 4016 982 4096 1016
rect 496 980 4096 982
rect 1674 970 1750 980
rect 1926 970 2002 980
rect 102 962 192 968
rect 408 856 442 872
rect 496 870 514 904
rect 548 870 582 904
rect 616 870 650 904
rect 684 870 718 904
rect 752 870 786 904
rect 820 870 854 904
rect 888 870 922 904
rect 956 870 990 904
rect 1024 870 1058 904
rect 1092 870 1126 904
rect 1160 870 1194 904
rect 1228 870 1262 904
rect 1296 870 1330 904
rect 1364 870 1398 904
rect 1432 870 1466 904
rect 1500 870 1804 904
rect 2374 900 2450 980
rect 408 806 442 822
rect 1598 752 1648 870
rect 1686 860 1804 870
rect 2370 898 2454 900
rect 2370 864 2396 898
rect 2430 864 2454 898
rect 2370 862 2454 864
rect 2676 878 4030 882
rect 1696 850 1804 860
rect 1710 838 1804 850
rect 1720 800 1804 838
rect 2244 816 2260 850
rect 2294 816 2310 850
rect 2676 844 2702 878
rect 2736 844 2866 878
rect 2900 844 3030 878
rect 3064 844 3194 878
rect 3228 844 3358 878
rect 3392 844 3522 878
rect 3556 844 3686 878
rect 3720 844 3764 878
rect 3798 844 3850 878
rect 3884 844 4030 878
rect 2676 840 4030 844
rect 1720 766 1746 800
rect 1780 766 1804 800
rect 2370 802 4132 804
rect 2370 774 2388 802
rect 2122 768 2388 774
rect 2422 768 4132 802
rect 1590 718 1606 752
rect 1640 718 1656 752
rect 260 698 1274 710
rect 260 664 314 698
rect 348 664 478 698
rect 512 664 642 698
rect 676 664 806 698
rect 840 664 970 698
rect 1004 664 1134 698
rect 1168 664 1274 698
rect 260 654 1274 664
rect 1720 670 1746 704
rect 1780 670 1804 704
rect 1720 654 1804 670
rect 2122 698 4132 768
rect 2122 696 2392 698
rect 2 620 42 654
rect 76 620 178 654
rect 212 620 314 654
rect 348 620 450 654
rect 484 620 586 654
rect 620 620 722 654
rect 756 620 858 654
rect 892 620 994 654
rect 1028 620 1130 654
rect 1164 620 1266 654
rect 1300 620 1402 654
rect 1436 620 1538 654
rect 1572 620 1674 654
rect 1708 620 1878 654
rect 1912 620 2014 654
rect 2048 620 2082 654
rect 186 460 224 620
rect 186 426 188 460
rect 222 426 224 460
rect 186 408 224 426
rect 282 542 334 552
rect 282 508 292 542
rect 326 508 334 542
rect 282 500 334 508
rect 282 460 320 500
rect 282 426 284 460
rect 318 426 320 460
rect 140 332 156 366
rect 190 332 206 366
rect 186 254 224 284
rect 186 220 188 254
rect 222 220 224 254
rect 186 182 224 220
rect 186 148 188 182
rect 222 148 224 182
rect 186 132 224 148
rect 282 276 320 426
rect 434 460 472 620
rect 802 546 1850 620
rect 2020 548 2054 564
rect 802 544 1884 546
rect 776 510 802 544
rect 836 510 932 544
rect 966 510 1000 544
rect 1034 510 1068 544
rect 1102 510 1136 544
rect 1170 510 1204 544
rect 1238 510 1272 544
rect 1306 510 1340 544
rect 1374 510 1408 544
rect 1442 510 1476 544
rect 1510 510 1544 544
rect 1578 510 1612 544
rect 1646 510 1680 544
rect 1714 510 1748 544
rect 1782 510 1816 544
rect 1850 510 1884 544
rect 924 508 1884 510
rect 2122 546 2192 696
rect 2228 620 2286 654
rect 2320 620 2422 654
rect 2456 620 2558 654
rect 2592 620 2694 654
rect 2728 620 2830 654
rect 2864 620 2966 654
rect 3000 620 3102 654
rect 3136 620 3238 654
rect 3272 620 3374 654
rect 3408 620 3510 654
rect 3544 620 3646 654
rect 3680 620 3782 654
rect 3816 620 3918 654
rect 3952 620 4132 654
rect 2416 608 3914 620
rect 2416 574 2470 608
rect 2504 574 2634 608
rect 2668 574 2798 608
rect 2832 574 2962 608
rect 2996 574 3126 608
rect 3160 574 3290 608
rect 3324 574 3446 608
rect 3480 574 3610 608
rect 3644 574 3774 608
rect 3808 574 3914 608
rect 2416 564 3914 574
rect 2020 498 2054 514
rect 2108 512 2140 546
rect 2174 512 2192 546
rect 434 426 436 460
rect 470 426 472 460
rect 434 408 472 426
rect 530 460 568 480
rect 530 426 532 460
rect 566 426 568 460
rect 388 332 404 366
rect 438 332 454 366
rect 530 348 568 426
rect 674 448 864 450
rect 674 414 690 448
rect 724 414 802 448
rect 836 414 864 448
rect 2108 444 2192 450
rect 1998 442 2192 444
rect 1998 434 2134 442
rect 674 412 864 414
rect 924 432 2134 434
rect 924 398 940 432
rect 974 398 1008 432
rect 1042 398 1076 432
rect 1110 398 1144 432
rect 1178 398 1212 432
rect 1246 398 1280 432
rect 1314 398 1348 432
rect 1382 398 1416 432
rect 1450 398 1484 432
rect 1518 398 1552 432
rect 1586 398 1620 432
rect 1654 398 1688 432
rect 1722 398 1756 432
rect 1790 398 1824 432
rect 1858 398 1892 432
rect 1926 408 2134 432
rect 2168 408 2192 442
rect 1926 398 2192 408
rect 924 396 2192 398
rect 530 329 862 348
rect 530 295 820 329
rect 854 295 862 329
rect 924 336 2230 338
rect 924 302 940 336
rect 974 302 1008 336
rect 1042 302 1076 336
rect 1110 302 1144 336
rect 1178 302 1212 336
rect 1246 302 1280 336
rect 1314 302 1348 336
rect 1382 302 1416 336
rect 1450 302 1484 336
rect 1518 302 1552 336
rect 1586 302 1620 336
rect 1654 302 1688 336
rect 1722 302 1756 336
rect 1790 302 1824 336
rect 1858 302 1892 336
rect 1926 302 2230 336
rect 924 300 2230 302
rect 282 242 284 276
rect 318 242 320 276
rect 282 208 320 242
rect 282 174 284 208
rect 318 174 320 208
rect 282 140 320 174
rect 434 256 472 284
rect 434 222 436 256
rect 470 222 472 256
rect 434 183 472 222
rect 434 148 436 183
rect 470 148 472 183
rect 434 132 472 148
rect 530 276 862 295
rect 530 242 532 276
rect 566 242 568 276
rect 530 208 568 242
rect 2034 220 2084 300
rect 2120 292 2230 300
rect 2134 284 2230 292
rect 2144 274 2230 284
rect 2146 268 2230 274
rect 2146 234 2172 268
rect 2206 234 2230 268
rect 530 174 532 208
rect 566 174 568 208
rect 2026 186 2042 220
rect 2076 186 2092 220
rect 530 140 568 174
rect 2146 178 2230 180
rect 644 134 780 146
rect 2146 138 2172 178
rect 2206 138 2230 178
rect 2320 156 2482 164
rect 644 100 686 134
rect 720 100 780 134
rect 644 64 780 100
rect 2320 122 2360 156
rect 2394 122 2482 156
rect 2320 64 2482 122
rect 0 30 42 64
rect 76 30 178 64
rect 212 30 314 64
rect 348 30 450 64
rect 484 30 586 64
rect 620 30 722 64
rect 756 30 858 64
rect 892 30 994 64
rect 1028 30 1130 64
rect 1164 30 1266 64
rect 1300 30 1402 64
rect 1436 30 1538 64
rect 1572 30 1674 64
rect 1708 30 1810 64
rect 1844 30 1946 64
rect 1980 30 2082 64
rect 2116 30 2218 64
rect 2252 30 2354 64
rect 2388 30 2490 64
rect 2524 30 2626 64
rect 2660 30 2762 64
rect 2796 30 2898 64
rect 2932 30 3034 64
rect 3068 30 3170 64
rect 3204 30 3306 64
rect 3340 30 3442 64
rect 3476 30 3578 64
rect 3612 30 3714 64
rect 3748 30 3850 64
rect 3884 30 3986 64
rect 4020 30 4134 64
<< viali >>
rect 42 1214 76 1248
rect 178 1214 212 1248
rect 314 1214 348 1248
rect 450 1214 484 1248
rect 586 1214 620 1248
rect 722 1214 756 1248
rect 858 1214 892 1248
rect 994 1214 1028 1248
rect 1130 1214 1164 1248
rect 1266 1214 1300 1248
rect 1402 1214 1436 1248
rect 1538 1214 1572 1248
rect 1674 1214 1708 1248
rect 1810 1214 1844 1248
rect 1946 1214 1980 1248
rect 2082 1214 2116 1248
rect 2218 1214 2252 1248
rect 2354 1214 2388 1248
rect 2490 1214 2524 1248
rect 2626 1214 2660 1248
rect 2762 1214 2796 1248
rect 2898 1214 2932 1248
rect 3034 1214 3068 1248
rect 3170 1214 3204 1248
rect 3306 1214 3340 1248
rect 3442 1214 3476 1248
rect 3578 1214 3612 1248
rect 3714 1214 3748 1248
rect 3850 1214 3884 1248
rect 3986 1214 4020 1248
rect 2562 1080 2588 1114
rect 2588 1080 2596 1114
rect 2646 1080 2656 1114
rect 2656 1080 2680 1114
rect 408 822 442 856
rect 2260 816 2294 850
rect 3764 844 3798 878
rect 3850 844 3884 878
rect 42 620 76 654
rect 178 620 212 654
rect 314 620 348 654
rect 450 620 484 654
rect 586 620 620 654
rect 722 620 756 654
rect 858 620 892 654
rect 994 620 1028 654
rect 1130 620 1164 654
rect 1266 620 1300 654
rect 1402 620 1436 654
rect 1538 620 1572 654
rect 1674 620 1708 654
rect 1878 620 1912 654
rect 2014 620 2048 654
rect 292 508 326 542
rect 156 332 190 366
rect 188 220 222 254
rect 188 148 222 182
rect 2020 514 2054 548
rect 2286 620 2320 654
rect 2422 620 2456 654
rect 2558 620 2592 654
rect 2694 620 2728 654
rect 2830 620 2864 654
rect 2966 620 3000 654
rect 3102 620 3136 654
rect 3238 620 3272 654
rect 3374 620 3408 654
rect 3510 620 3544 654
rect 3646 620 3680 654
rect 3782 620 3816 654
rect 3918 620 3952 654
rect 404 332 438 366
rect 436 222 470 256
rect 436 182 470 183
rect 436 149 470 182
rect 2172 172 2206 178
rect 2172 144 2206 172
rect 42 30 76 64
rect 178 30 212 64
rect 314 30 348 64
rect 450 30 484 64
rect 586 30 620 64
rect 722 30 756 64
rect 858 30 892 64
rect 994 30 1028 64
rect 1130 30 1164 64
rect 1266 30 1300 64
rect 1402 30 1436 64
rect 1538 30 1572 64
rect 1674 30 1708 64
rect 1810 30 1844 64
rect 1946 30 1980 64
rect 2082 30 2116 64
rect 2218 30 2252 64
rect 2354 30 2388 64
rect 2490 30 2524 64
rect 2626 30 2660 64
rect 2762 30 2796 64
rect 2898 30 2932 64
rect 3034 30 3068 64
rect 3170 30 3204 64
rect 3306 30 3340 64
rect 3442 30 3476 64
rect 3578 30 3612 64
rect 3714 30 3748 64
rect 3850 30 3884 64
rect 3986 30 4020 64
<< metal1 >>
rect 0 1248 4132 1280
rect 0 1214 42 1248
rect 76 1214 178 1248
rect 212 1214 314 1248
rect 348 1214 450 1248
rect 484 1214 586 1248
rect 620 1214 722 1248
rect 756 1214 858 1248
rect 892 1214 994 1248
rect 1028 1214 1130 1248
rect 1164 1214 1266 1248
rect 1300 1214 1402 1248
rect 1436 1214 1538 1248
rect 1572 1214 1674 1248
rect 1708 1214 1810 1248
rect 1844 1214 1946 1248
rect 1980 1214 2082 1248
rect 2116 1214 2218 1248
rect 2252 1214 2354 1248
rect 2388 1214 2490 1248
rect 2524 1214 2626 1248
rect 2660 1214 2762 1248
rect 2796 1214 2898 1248
rect 2932 1214 3034 1248
rect 3068 1214 3170 1248
rect 3204 1214 3306 1248
rect 3340 1214 3442 1248
rect 3476 1214 3578 1248
rect 3612 1214 3714 1248
rect 3748 1214 3850 1248
rect 3884 1214 3986 1248
rect 4020 1214 4132 1248
rect 0 1184 4132 1214
rect 2550 1120 2686 1126
rect 2550 1114 2586 1120
rect 2638 1114 2686 1120
rect 2550 1080 2562 1114
rect 2638 1080 2646 1114
rect 2680 1080 2686 1114
rect 2550 1068 2586 1080
rect 2638 1068 2686 1080
rect 3752 892 3892 1184
rect 3752 878 3896 892
rect 392 864 456 870
rect 392 812 398 864
rect 450 812 456 864
rect 392 806 456 812
rect 2244 858 2308 864
rect 2244 806 2250 858
rect 2302 806 2308 858
rect 3752 844 3764 878
rect 3798 844 3850 878
rect 3884 844 3896 878
rect 3752 832 3896 844
rect 2244 804 2308 806
rect 2 654 4132 688
rect 2 620 42 654
rect 76 620 178 654
rect 212 620 314 654
rect 348 620 450 654
rect 484 620 586 654
rect 620 620 722 654
rect 756 620 858 654
rect 892 620 994 654
rect 1028 620 1130 654
rect 1164 620 1266 654
rect 1300 620 1402 654
rect 1436 620 1538 654
rect 1572 620 1674 654
rect 1708 620 1878 654
rect 1912 620 2014 654
rect 2048 620 2286 654
rect 2320 620 2422 654
rect 2456 620 2558 654
rect 2592 620 2694 654
rect 2728 620 2830 654
rect 2864 620 2966 654
rect 3000 620 3102 654
rect 3136 620 3238 654
rect 3272 620 3374 654
rect 3408 620 3510 654
rect 3544 620 3646 654
rect 3680 620 3782 654
rect 3816 620 3918 654
rect 3952 620 4132 654
rect 2 592 4132 620
rect 2004 556 2068 562
rect 276 550 340 556
rect 276 498 282 550
rect 334 498 340 550
rect 2004 504 2010 556
rect 2062 504 2068 556
rect 2004 498 2068 504
rect 276 492 340 498
rect 2536 410 2694 458
rect 142 374 206 380
rect 142 322 148 374
rect 200 322 206 374
rect 142 316 206 322
rect 388 374 452 380
rect 388 322 394 374
rect 446 322 452 374
rect 388 316 452 322
rect 2536 358 2590 410
rect 2642 358 2694 410
rect 2536 308 2694 358
rect 180 254 230 266
rect 180 220 188 254
rect 222 220 230 254
rect 180 198 230 220
rect 428 256 478 268
rect 428 222 436 256
rect 470 222 478 256
rect 428 198 478 222
rect 2536 198 2632 308
rect 180 183 2632 198
rect 180 182 436 183
rect 180 148 188 182
rect 222 149 436 182
rect 470 178 2632 183
rect 470 149 2172 178
rect 222 148 2172 149
rect 180 144 2172 148
rect 2206 144 2632 178
rect 180 138 2632 144
rect 180 136 226 138
rect 436 130 470 138
rect 0 64 4134 96
rect 0 30 42 64
rect 76 30 178 64
rect 212 30 314 64
rect 348 30 450 64
rect 484 30 586 64
rect 620 30 722 64
rect 756 30 858 64
rect 892 30 994 64
rect 1028 30 1130 64
rect 1164 30 1266 64
rect 1300 30 1402 64
rect 1436 30 1538 64
rect 1572 30 1674 64
rect 1708 30 1810 64
rect 1844 30 1946 64
rect 1980 30 2082 64
rect 2116 30 2218 64
rect 2252 30 2354 64
rect 2388 30 2490 64
rect 2524 30 2626 64
rect 2660 30 2762 64
rect 2796 30 2898 64
rect 2932 30 3034 64
rect 3068 30 3170 64
rect 3204 30 3306 64
rect 3340 30 3442 64
rect 3476 30 3578 64
rect 3612 30 3714 64
rect 3748 30 3850 64
rect 3884 30 3986 64
rect 4020 30 4134 64
rect 0 0 4134 30
<< via1 >>
rect 2586 1114 2638 1120
rect 2586 1080 2596 1114
rect 2596 1080 2638 1114
rect 2586 1068 2638 1080
rect 398 856 450 864
rect 398 822 408 856
rect 408 822 442 856
rect 442 822 450 856
rect 398 812 450 822
rect 2250 850 2302 858
rect 2250 816 2260 850
rect 2260 816 2294 850
rect 2294 816 2302 850
rect 2250 806 2302 816
rect 282 542 334 550
rect 282 508 292 542
rect 292 508 326 542
rect 326 508 334 542
rect 282 498 334 508
rect 2010 548 2062 556
rect 2010 514 2020 548
rect 2020 514 2054 548
rect 2054 514 2062 548
rect 2010 504 2062 514
rect 148 366 200 374
rect 148 332 156 366
rect 156 332 190 366
rect 190 332 200 366
rect 148 322 200 332
rect 394 366 446 374
rect 394 332 404 366
rect 404 332 438 366
rect 438 332 446 366
rect 394 322 446 332
rect 2590 358 2642 410
<< metal2 >>
rect 2556 1120 2678 1126
rect 2556 1068 2586 1120
rect 2638 1068 2678 1120
rect 368 866 456 870
rect 120 864 456 866
rect 120 812 398 864
rect 450 812 456 864
rect 120 806 456 812
rect 1740 858 2308 864
rect 1740 806 2250 858
rect 2302 806 2308 858
rect 120 794 454 806
rect 1740 800 2308 806
rect 120 544 184 794
rect 1740 600 1834 800
rect 2 482 184 544
rect 276 550 1834 600
rect 276 498 282 550
rect 334 520 1834 550
rect 1894 556 2068 562
rect 334 498 340 520
rect 276 492 340 498
rect 1894 504 2010 556
rect 2062 504 2068 556
rect 1894 498 2068 504
rect 120 380 184 482
rect 120 374 206 380
rect 120 322 148 374
rect 200 322 206 374
rect 120 316 206 322
rect 352 374 452 380
rect 352 322 394 374
rect 446 322 452 374
rect 352 220 418 322
rect 1894 220 1968 498
rect 2556 410 2678 1068
rect 2556 358 2590 410
rect 2642 358 2678 410
rect 2556 342 2678 358
rect 352 218 1968 220
rect 2 146 1968 218
<< labels >>
rlabel metal1 s 0 48 0 48 4 VDD
port 1 nsew
rlabel metal1 s 0 1232 0 1232 4 VDD
port 1 nsew
rlabel metal1 s 2 640 2 640 4 GND
port 2 nsew
rlabel metal2 s 2 182 2 182 4 Up
port 3 nsew
rlabel metal2 s 2 512 2 512 4 Down
port 4 nsew
rlabel locali s 4132 750 4132 750 4 Out
port 5 nsew
rlabel locali s 102 986 102 986 4 ENb
port 6 nsew
<< end >>
