* SPICE3 file created from dram_cell.ext - technology: sky130A

.subckt dram_cell WWL WBL RWL RBL
X0 RWL a_50_n70# RBL VSUBS sky130_fd_pr__nfet_01v8 ad=3e+11p pd=2.6e+06u as=3.5e+11p ps=2.7e+06u w=1e+06u l=150000u
X1 a_50_n70# WWL WBL VSUBS sky130_fd_pr__nfet_01v8 ad=3.5e+11p pd=2.7e+06u as=3e+11p ps=2.6e+06u w=1e+06u l=150000u
.ends

