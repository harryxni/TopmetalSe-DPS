magic
tech sky130B
magscale 1 2
timestamp 1661296583
<< poly >>
rect 60 -65 90 30
rect 60 -323 90 -280
rect 7 -333 90 -323
rect 7 -367 23 -333
rect 57 -365 90 -333
rect 57 -367 73 -365
rect 7 -377 73 -367
<< polycont >>
rect 23 -367 57 -333
<< locali >>
rect 0 210 40 270
rect 350 197 380 230
rect 350 115 380 163
rect 230 20 253 50
rect 0 -120 40 -80
rect 0 -280 40 -260
rect 23 -333 57 -317
rect 23 -383 57 -367
<< viali >>
rect 0 270 40 310
rect 348 163 382 197
rect 253 18 287 52
rect 228 -102 262 -68
rect 0 -160 40 -120
rect 23 -367 57 -333
<< metal1 >>
rect -6 316 46 322
rect -12 264 -6 316
rect 46 264 52 316
rect -6 258 46 264
rect 342 206 388 209
rect 333 154 339 206
rect 391 154 397 206
rect 342 151 388 154
rect 244 61 296 67
rect 244 3 296 9
rect 219 -59 271 -53
rect -10 -114 50 -100
rect 216 -108 219 -62
rect -12 -120 50 -114
rect 271 -108 274 -62
rect 219 -117 271 -111
rect -12 -160 0 -120
rect 40 -160 50 -120
rect -12 -166 50 -160
rect -10 -180 50 -166
rect 78 -180 84 -174
rect -10 -220 84 -180
rect 78 -226 84 -220
rect 136 -226 142 -174
rect 17 -333 63 -321
rect 268 -333 274 -324
rect 17 -367 23 -333
rect 57 -367 274 -333
rect 17 -379 63 -367
rect 268 -376 274 -367
rect 326 -376 332 -324
<< via1 >>
rect -6 310 46 316
rect -6 270 0 310
rect 0 270 40 310
rect 40 270 46 310
rect -6 264 46 270
rect 339 197 391 206
rect 339 163 348 197
rect 348 163 382 197
rect 382 163 391 197
rect 339 154 391 163
rect 244 52 296 61
rect 244 18 253 52
rect 253 18 287 52
rect 287 18 296 52
rect 244 9 296 18
rect 219 -68 271 -59
rect 219 -102 228 -68
rect 228 -102 262 -68
rect 262 -102 271 -68
rect 219 -111 271 -102
rect 84 -226 136 -174
rect 274 -376 326 -324
<< metal2 >>
rect 0 316 40 370
rect -12 264 -6 316
rect 46 264 52 316
rect 0 -430 40 264
rect 175 -50 205 370
rect 339 210 391 212
rect 326 150 335 210
rect 395 150 404 210
rect 339 148 391 150
rect 261 61 270 65
rect 238 9 244 61
rect 261 5 270 9
rect 330 5 339 65
rect 175 -59 280 -50
rect 175 -111 219 -59
rect 271 -111 280 -59
rect 175 -120 280 -111
rect 70 -170 140 -160
rect 70 -230 80 -170
rect 70 -240 140 -230
rect 175 -430 205 -120
rect 274 -320 326 -318
rect 261 -380 270 -320
rect 330 -380 339 -320
rect 274 -382 326 -380
<< via2 >>
rect 335 206 395 210
rect 335 154 339 206
rect 339 154 391 206
rect 391 154 395 206
rect 335 150 395 154
rect 270 61 330 65
rect 270 9 296 61
rect 296 9 330 61
rect 270 5 330 9
rect 80 -174 140 -170
rect 80 -226 84 -174
rect 84 -226 136 -174
rect 136 -226 140 -174
rect 80 -230 140 -226
rect 270 -324 330 -320
rect 270 -376 274 -324
rect 274 -376 326 -324
rect 326 -376 330 -324
rect 270 -380 330 -376
<< metal3 >>
rect 330 210 400 215
rect -60 150 335 210
rect 395 150 420 210
rect 330 145 400 150
rect 265 70 335 76
rect 240 6 265 70
rect 335 6 340 70
rect 240 5 270 6
rect 330 5 340 6
rect 240 0 340 5
rect 265 -50 335 0
rect 60 -165 160 -120
rect 60 -235 75 -165
rect 145 -235 160 -165
rect 60 -260 160 -235
rect 265 -320 335 -315
rect -90 -380 270 -320
rect 330 -380 420 -320
rect 265 -385 335 -380
<< via3 >>
rect 265 65 335 70
rect 265 6 270 65
rect 270 6 330 65
rect 330 6 335 65
rect 75 -170 145 -165
rect 75 -230 80 -170
rect 80 -230 140 -170
rect 140 -230 145 -170
rect 75 -235 145 -230
<< metal4 >>
rect 80 -164 140 370
rect 270 71 330 370
rect 264 70 336 71
rect 264 6 265 70
rect 335 6 336 70
rect 264 5 336 6
rect 74 -165 146 -164
rect 74 -235 75 -165
rect 145 -235 146 -165
rect 74 -236 146 -235
rect 80 -430 140 -236
rect 270 -430 330 5
use dram_cell  dram_cell_0
timestamp 1660883971
transform 1 0 40 0 1 100
box -40 -100 340 223
use dram_cell  dram_cell_1
timestamp 1660883971
transform 1 0 40 0 -1 -150
box -40 -100 340 223
<< labels >>
rlabel space 60 -340 90 55 3 TEST
port 8 e
rlabel space 60 -375 90 30 3 test
<< end >>
