magic
tech sky130B
magscale 1 2
timestamp 1606426375
<< error_p >>
rect -1740 381 -1682 387
rect -1622 381 -1564 387
rect -1504 381 -1446 387
rect -1386 381 -1328 387
rect -1268 381 -1210 387
rect -1150 381 -1092 387
rect -1032 381 -974 387
rect -914 381 -856 387
rect -796 381 -738 387
rect -678 381 -620 387
rect -560 381 -502 387
rect -442 381 -384 387
rect -324 381 -266 387
rect -206 381 -148 387
rect -88 381 -30 387
rect 30 381 88 387
rect 148 381 206 387
rect 266 381 324 387
rect 384 381 442 387
rect 502 381 560 387
rect 620 381 678 387
rect 738 381 796 387
rect 856 381 914 387
rect 974 381 1032 387
rect 1092 381 1150 387
rect 1210 381 1268 387
rect 1328 381 1386 387
rect 1446 381 1504 387
rect 1564 381 1622 387
rect 1682 381 1740 387
rect -1740 347 -1728 381
rect -1622 347 -1610 381
rect -1504 347 -1492 381
rect -1386 347 -1374 381
rect -1268 347 -1256 381
rect -1150 347 -1138 381
rect -1032 347 -1020 381
rect -914 347 -902 381
rect -796 347 -784 381
rect -678 347 -666 381
rect -560 347 -548 381
rect -442 347 -430 381
rect -324 347 -312 381
rect -206 347 -194 381
rect -88 347 -76 381
rect 30 347 42 381
rect 148 347 160 381
rect 266 347 278 381
rect 384 347 396 381
rect 502 347 514 381
rect 620 347 632 381
rect 738 347 750 381
rect 856 347 868 381
rect 974 347 986 381
rect 1092 347 1104 381
rect 1210 347 1222 381
rect 1328 347 1340 381
rect 1446 347 1458 381
rect 1564 347 1576 381
rect 1682 347 1694 381
rect -1740 341 -1682 347
rect -1622 341 -1564 347
rect -1504 341 -1446 347
rect -1386 341 -1328 347
rect -1268 341 -1210 347
rect -1150 341 -1092 347
rect -1032 341 -974 347
rect -914 341 -856 347
rect -796 341 -738 347
rect -678 341 -620 347
rect -560 341 -502 347
rect -442 341 -384 347
rect -324 341 -266 347
rect -206 341 -148 347
rect -88 341 -30 347
rect 30 341 88 347
rect 148 341 206 347
rect 266 341 324 347
rect 384 341 442 347
rect 502 341 560 347
rect 620 341 678 347
rect 738 341 796 347
rect 856 341 914 347
rect 974 341 1032 347
rect 1092 341 1150 347
rect 1210 341 1268 347
rect 1328 341 1386 347
rect 1446 341 1504 347
rect 1564 341 1622 347
rect 1682 341 1740 347
rect -1740 -347 -1682 -341
rect -1622 -347 -1564 -341
rect -1504 -347 -1446 -341
rect -1386 -347 -1328 -341
rect -1268 -347 -1210 -341
rect -1150 -347 -1092 -341
rect -1032 -347 -974 -341
rect -914 -347 -856 -341
rect -796 -347 -738 -341
rect -678 -347 -620 -341
rect -560 -347 -502 -341
rect -442 -347 -384 -341
rect -324 -347 -266 -341
rect -206 -347 -148 -341
rect -88 -347 -30 -341
rect 30 -347 88 -341
rect 148 -347 206 -341
rect 266 -347 324 -341
rect 384 -347 442 -341
rect 502 -347 560 -341
rect 620 -347 678 -341
rect 738 -347 796 -341
rect 856 -347 914 -341
rect 974 -347 1032 -341
rect 1092 -347 1150 -341
rect 1210 -347 1268 -341
rect 1328 -347 1386 -341
rect 1446 -347 1504 -341
rect 1564 -347 1622 -341
rect 1682 -347 1740 -341
rect -1740 -381 -1728 -347
rect -1622 -381 -1610 -347
rect -1504 -381 -1492 -347
rect -1386 -381 -1374 -347
rect -1268 -381 -1256 -347
rect -1150 -381 -1138 -347
rect -1032 -381 -1020 -347
rect -914 -381 -902 -347
rect -796 -381 -784 -347
rect -678 -381 -666 -347
rect -560 -381 -548 -347
rect -442 -381 -430 -347
rect -324 -381 -312 -347
rect -206 -381 -194 -347
rect -88 -381 -76 -347
rect 30 -381 42 -347
rect 148 -381 160 -347
rect 266 -381 278 -347
rect 384 -381 396 -347
rect 502 -381 514 -347
rect 620 -381 632 -347
rect 738 -381 750 -347
rect 856 -381 868 -347
rect 974 -381 986 -347
rect 1092 -381 1104 -347
rect 1210 -381 1222 -347
rect 1328 -381 1340 -347
rect 1446 -381 1458 -347
rect 1564 -381 1576 -347
rect 1682 -381 1694 -347
rect -1740 -387 -1682 -381
rect -1622 -387 -1564 -381
rect -1504 -387 -1446 -381
rect -1386 -387 -1328 -381
rect -1268 -387 -1210 -381
rect -1150 -387 -1092 -381
rect -1032 -387 -974 -381
rect -914 -387 -856 -381
rect -796 -387 -738 -381
rect -678 -387 -620 -381
rect -560 -387 -502 -381
rect -442 -387 -384 -381
rect -324 -387 -266 -381
rect -206 -387 -148 -381
rect -88 -387 -30 -381
rect 30 -387 88 -381
rect 148 -387 206 -381
rect 266 -387 324 -381
rect 384 -387 442 -381
rect 502 -387 560 -381
rect 620 -387 678 -381
rect 738 -387 796 -381
rect 856 -387 914 -381
rect 974 -387 1032 -381
rect 1092 -387 1150 -381
rect 1210 -387 1268 -381
rect 1328 -387 1386 -381
rect 1446 -387 1504 -381
rect 1564 -387 1622 -381
rect 1682 -387 1740 -381
<< nwell >>
rect -1937 -519 1937 519
<< pmos >>
rect -1741 -300 -1681 300
rect -1623 -300 -1563 300
rect -1505 -300 -1445 300
rect -1387 -300 -1327 300
rect -1269 -300 -1209 300
rect -1151 -300 -1091 300
rect -1033 -300 -973 300
rect -915 -300 -855 300
rect -797 -300 -737 300
rect -679 -300 -619 300
rect -561 -300 -501 300
rect -443 -300 -383 300
rect -325 -300 -265 300
rect -207 -300 -147 300
rect -89 -300 -29 300
rect 29 -300 89 300
rect 147 -300 207 300
rect 265 -300 325 300
rect 383 -300 443 300
rect 501 -300 561 300
rect 619 -300 679 300
rect 737 -300 797 300
rect 855 -300 915 300
rect 973 -300 1033 300
rect 1091 -300 1151 300
rect 1209 -300 1269 300
rect 1327 -300 1387 300
rect 1445 -300 1505 300
rect 1563 -300 1623 300
rect 1681 -300 1741 300
<< pdiff >>
rect -1799 288 -1741 300
rect -1799 -288 -1787 288
rect -1753 -288 -1741 288
rect -1799 -300 -1741 -288
rect -1681 288 -1623 300
rect -1681 -288 -1669 288
rect -1635 -288 -1623 288
rect -1681 -300 -1623 -288
rect -1563 288 -1505 300
rect -1563 -288 -1551 288
rect -1517 -288 -1505 288
rect -1563 -300 -1505 -288
rect -1445 288 -1387 300
rect -1445 -288 -1433 288
rect -1399 -288 -1387 288
rect -1445 -300 -1387 -288
rect -1327 288 -1269 300
rect -1327 -288 -1315 288
rect -1281 -288 -1269 288
rect -1327 -300 -1269 -288
rect -1209 288 -1151 300
rect -1209 -288 -1197 288
rect -1163 -288 -1151 288
rect -1209 -300 -1151 -288
rect -1091 288 -1033 300
rect -1091 -288 -1079 288
rect -1045 -288 -1033 288
rect -1091 -300 -1033 -288
rect -973 288 -915 300
rect -973 -288 -961 288
rect -927 -288 -915 288
rect -973 -300 -915 -288
rect -855 288 -797 300
rect -855 -288 -843 288
rect -809 -288 -797 288
rect -855 -300 -797 -288
rect -737 288 -679 300
rect -737 -288 -725 288
rect -691 -288 -679 288
rect -737 -300 -679 -288
rect -619 288 -561 300
rect -619 -288 -607 288
rect -573 -288 -561 288
rect -619 -300 -561 -288
rect -501 288 -443 300
rect -501 -288 -489 288
rect -455 -288 -443 288
rect -501 -300 -443 -288
rect -383 288 -325 300
rect -383 -288 -371 288
rect -337 -288 -325 288
rect -383 -300 -325 -288
rect -265 288 -207 300
rect -265 -288 -253 288
rect -219 -288 -207 288
rect -265 -300 -207 -288
rect -147 288 -89 300
rect -147 -288 -135 288
rect -101 -288 -89 288
rect -147 -300 -89 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 89 288 147 300
rect 89 -288 101 288
rect 135 -288 147 288
rect 89 -300 147 -288
rect 207 288 265 300
rect 207 -288 219 288
rect 253 -288 265 288
rect 207 -300 265 -288
rect 325 288 383 300
rect 325 -288 337 288
rect 371 -288 383 288
rect 325 -300 383 -288
rect 443 288 501 300
rect 443 -288 455 288
rect 489 -288 501 288
rect 443 -300 501 -288
rect 561 288 619 300
rect 561 -288 573 288
rect 607 -288 619 288
rect 561 -300 619 -288
rect 679 288 737 300
rect 679 -288 691 288
rect 725 -288 737 288
rect 679 -300 737 -288
rect 797 288 855 300
rect 797 -288 809 288
rect 843 -288 855 288
rect 797 -300 855 -288
rect 915 288 973 300
rect 915 -288 927 288
rect 961 -288 973 288
rect 915 -300 973 -288
rect 1033 288 1091 300
rect 1033 -288 1045 288
rect 1079 -288 1091 288
rect 1033 -300 1091 -288
rect 1151 288 1209 300
rect 1151 -288 1163 288
rect 1197 -288 1209 288
rect 1151 -300 1209 -288
rect 1269 288 1327 300
rect 1269 -288 1281 288
rect 1315 -288 1327 288
rect 1269 -300 1327 -288
rect 1387 288 1445 300
rect 1387 -288 1399 288
rect 1433 -288 1445 288
rect 1387 -300 1445 -288
rect 1505 288 1563 300
rect 1505 -288 1517 288
rect 1551 -288 1563 288
rect 1505 -300 1563 -288
rect 1623 288 1681 300
rect 1623 -288 1635 288
rect 1669 -288 1681 288
rect 1623 -300 1681 -288
rect 1741 288 1799 300
rect 1741 -288 1753 288
rect 1787 -288 1799 288
rect 1741 -300 1799 -288
<< pdiffc >>
rect -1787 -288 -1753 288
rect -1669 -288 -1635 288
rect -1551 -288 -1517 288
rect -1433 -288 -1399 288
rect -1315 -288 -1281 288
rect -1197 -288 -1163 288
rect -1079 -288 -1045 288
rect -961 -288 -927 288
rect -843 -288 -809 288
rect -725 -288 -691 288
rect -607 -288 -573 288
rect -489 -288 -455 288
rect -371 -288 -337 288
rect -253 -288 -219 288
rect -135 -288 -101 288
rect -17 -288 17 288
rect 101 -288 135 288
rect 219 -288 253 288
rect 337 -288 371 288
rect 455 -288 489 288
rect 573 -288 607 288
rect 691 -288 725 288
rect 809 -288 843 288
rect 927 -288 961 288
rect 1045 -288 1079 288
rect 1163 -288 1197 288
rect 1281 -288 1315 288
rect 1399 -288 1433 288
rect 1517 -288 1551 288
rect 1635 -288 1669 288
rect 1753 -288 1787 288
<< nsubdiff >>
rect -1901 449 -1805 483
rect 1805 449 1901 483
rect -1901 387 -1867 449
rect 1867 387 1901 449
rect -1901 -449 -1867 -387
rect 1867 -449 1901 -387
rect -1901 -483 -1805 -449
rect 1805 -483 1901 -449
<< nsubdiffcont >>
rect -1805 449 1805 483
rect -1901 -387 -1867 387
rect 1867 -387 1901 387
rect -1805 -483 1805 -449
<< poly >>
rect -1744 381 -1678 397
rect -1744 347 -1728 381
rect -1694 347 -1678 381
rect -1744 331 -1678 347
rect -1626 381 -1560 397
rect -1626 347 -1610 381
rect -1576 347 -1560 381
rect -1626 331 -1560 347
rect -1508 381 -1442 397
rect -1508 347 -1492 381
rect -1458 347 -1442 381
rect -1508 331 -1442 347
rect -1390 381 -1324 397
rect -1390 347 -1374 381
rect -1340 347 -1324 381
rect -1390 331 -1324 347
rect -1272 381 -1206 397
rect -1272 347 -1256 381
rect -1222 347 -1206 381
rect -1272 331 -1206 347
rect -1154 381 -1088 397
rect -1154 347 -1138 381
rect -1104 347 -1088 381
rect -1154 331 -1088 347
rect -1036 381 -970 397
rect -1036 347 -1020 381
rect -986 347 -970 381
rect -1036 331 -970 347
rect -918 381 -852 397
rect -918 347 -902 381
rect -868 347 -852 381
rect -918 331 -852 347
rect -800 381 -734 397
rect -800 347 -784 381
rect -750 347 -734 381
rect -800 331 -734 347
rect -682 381 -616 397
rect -682 347 -666 381
rect -632 347 -616 381
rect -682 331 -616 347
rect -564 381 -498 397
rect -564 347 -548 381
rect -514 347 -498 381
rect -564 331 -498 347
rect -446 381 -380 397
rect -446 347 -430 381
rect -396 347 -380 381
rect -446 331 -380 347
rect -328 381 -262 397
rect -328 347 -312 381
rect -278 347 -262 381
rect -328 331 -262 347
rect -210 381 -144 397
rect -210 347 -194 381
rect -160 347 -144 381
rect -210 331 -144 347
rect -92 381 -26 397
rect -92 347 -76 381
rect -42 347 -26 381
rect -92 331 -26 347
rect 26 381 92 397
rect 26 347 42 381
rect 76 347 92 381
rect 26 331 92 347
rect 144 381 210 397
rect 144 347 160 381
rect 194 347 210 381
rect 144 331 210 347
rect 262 381 328 397
rect 262 347 278 381
rect 312 347 328 381
rect 262 331 328 347
rect 380 381 446 397
rect 380 347 396 381
rect 430 347 446 381
rect 380 331 446 347
rect 498 381 564 397
rect 498 347 514 381
rect 548 347 564 381
rect 498 331 564 347
rect 616 381 682 397
rect 616 347 632 381
rect 666 347 682 381
rect 616 331 682 347
rect 734 381 800 397
rect 734 347 750 381
rect 784 347 800 381
rect 734 331 800 347
rect 852 381 918 397
rect 852 347 868 381
rect 902 347 918 381
rect 852 331 918 347
rect 970 381 1036 397
rect 970 347 986 381
rect 1020 347 1036 381
rect 970 331 1036 347
rect 1088 381 1154 397
rect 1088 347 1104 381
rect 1138 347 1154 381
rect 1088 331 1154 347
rect 1206 381 1272 397
rect 1206 347 1222 381
rect 1256 347 1272 381
rect 1206 331 1272 347
rect 1324 381 1390 397
rect 1324 347 1340 381
rect 1374 347 1390 381
rect 1324 331 1390 347
rect 1442 381 1508 397
rect 1442 347 1458 381
rect 1492 347 1508 381
rect 1442 331 1508 347
rect 1560 381 1626 397
rect 1560 347 1576 381
rect 1610 347 1626 381
rect 1560 331 1626 347
rect 1678 381 1744 397
rect 1678 347 1694 381
rect 1728 347 1744 381
rect 1678 331 1744 347
rect -1741 300 -1681 331
rect -1623 300 -1563 331
rect -1505 300 -1445 331
rect -1387 300 -1327 331
rect -1269 300 -1209 331
rect -1151 300 -1091 331
rect -1033 300 -973 331
rect -915 300 -855 331
rect -797 300 -737 331
rect -679 300 -619 331
rect -561 300 -501 331
rect -443 300 -383 331
rect -325 300 -265 331
rect -207 300 -147 331
rect -89 300 -29 331
rect 29 300 89 331
rect 147 300 207 331
rect 265 300 325 331
rect 383 300 443 331
rect 501 300 561 331
rect 619 300 679 331
rect 737 300 797 331
rect 855 300 915 331
rect 973 300 1033 331
rect 1091 300 1151 331
rect 1209 300 1269 331
rect 1327 300 1387 331
rect 1445 300 1505 331
rect 1563 300 1623 331
rect 1681 300 1741 331
rect -1741 -331 -1681 -300
rect -1623 -331 -1563 -300
rect -1505 -331 -1445 -300
rect -1387 -331 -1327 -300
rect -1269 -331 -1209 -300
rect -1151 -331 -1091 -300
rect -1033 -331 -973 -300
rect -915 -331 -855 -300
rect -797 -331 -737 -300
rect -679 -331 -619 -300
rect -561 -331 -501 -300
rect -443 -331 -383 -300
rect -325 -331 -265 -300
rect -207 -331 -147 -300
rect -89 -331 -29 -300
rect 29 -331 89 -300
rect 147 -331 207 -300
rect 265 -331 325 -300
rect 383 -331 443 -300
rect 501 -331 561 -300
rect 619 -331 679 -300
rect 737 -331 797 -300
rect 855 -331 915 -300
rect 973 -331 1033 -300
rect 1091 -331 1151 -300
rect 1209 -331 1269 -300
rect 1327 -331 1387 -300
rect 1445 -331 1505 -300
rect 1563 -331 1623 -300
rect 1681 -331 1741 -300
rect -1744 -347 -1678 -331
rect -1744 -381 -1728 -347
rect -1694 -381 -1678 -347
rect -1744 -397 -1678 -381
rect -1626 -347 -1560 -331
rect -1626 -381 -1610 -347
rect -1576 -381 -1560 -347
rect -1626 -397 -1560 -381
rect -1508 -347 -1442 -331
rect -1508 -381 -1492 -347
rect -1458 -381 -1442 -347
rect -1508 -397 -1442 -381
rect -1390 -347 -1324 -331
rect -1390 -381 -1374 -347
rect -1340 -381 -1324 -347
rect -1390 -397 -1324 -381
rect -1272 -347 -1206 -331
rect -1272 -381 -1256 -347
rect -1222 -381 -1206 -347
rect -1272 -397 -1206 -381
rect -1154 -347 -1088 -331
rect -1154 -381 -1138 -347
rect -1104 -381 -1088 -347
rect -1154 -397 -1088 -381
rect -1036 -347 -970 -331
rect -1036 -381 -1020 -347
rect -986 -381 -970 -347
rect -1036 -397 -970 -381
rect -918 -347 -852 -331
rect -918 -381 -902 -347
rect -868 -381 -852 -347
rect -918 -397 -852 -381
rect -800 -347 -734 -331
rect -800 -381 -784 -347
rect -750 -381 -734 -347
rect -800 -397 -734 -381
rect -682 -347 -616 -331
rect -682 -381 -666 -347
rect -632 -381 -616 -347
rect -682 -397 -616 -381
rect -564 -347 -498 -331
rect -564 -381 -548 -347
rect -514 -381 -498 -347
rect -564 -397 -498 -381
rect -446 -347 -380 -331
rect -446 -381 -430 -347
rect -396 -381 -380 -347
rect -446 -397 -380 -381
rect -328 -347 -262 -331
rect -328 -381 -312 -347
rect -278 -381 -262 -347
rect -328 -397 -262 -381
rect -210 -347 -144 -331
rect -210 -381 -194 -347
rect -160 -381 -144 -347
rect -210 -397 -144 -381
rect -92 -347 -26 -331
rect -92 -381 -76 -347
rect -42 -381 -26 -347
rect -92 -397 -26 -381
rect 26 -347 92 -331
rect 26 -381 42 -347
rect 76 -381 92 -347
rect 26 -397 92 -381
rect 144 -347 210 -331
rect 144 -381 160 -347
rect 194 -381 210 -347
rect 144 -397 210 -381
rect 262 -347 328 -331
rect 262 -381 278 -347
rect 312 -381 328 -347
rect 262 -397 328 -381
rect 380 -347 446 -331
rect 380 -381 396 -347
rect 430 -381 446 -347
rect 380 -397 446 -381
rect 498 -347 564 -331
rect 498 -381 514 -347
rect 548 -381 564 -347
rect 498 -397 564 -381
rect 616 -347 682 -331
rect 616 -381 632 -347
rect 666 -381 682 -347
rect 616 -397 682 -381
rect 734 -347 800 -331
rect 734 -381 750 -347
rect 784 -381 800 -347
rect 734 -397 800 -381
rect 852 -347 918 -331
rect 852 -381 868 -347
rect 902 -381 918 -347
rect 852 -397 918 -381
rect 970 -347 1036 -331
rect 970 -381 986 -347
rect 1020 -381 1036 -347
rect 970 -397 1036 -381
rect 1088 -347 1154 -331
rect 1088 -381 1104 -347
rect 1138 -381 1154 -347
rect 1088 -397 1154 -381
rect 1206 -347 1272 -331
rect 1206 -381 1222 -347
rect 1256 -381 1272 -347
rect 1206 -397 1272 -381
rect 1324 -347 1390 -331
rect 1324 -381 1340 -347
rect 1374 -381 1390 -347
rect 1324 -397 1390 -381
rect 1442 -347 1508 -331
rect 1442 -381 1458 -347
rect 1492 -381 1508 -347
rect 1442 -397 1508 -381
rect 1560 -347 1626 -331
rect 1560 -381 1576 -347
rect 1610 -381 1626 -347
rect 1560 -397 1626 -381
rect 1678 -347 1744 -331
rect 1678 -381 1694 -347
rect 1728 -381 1744 -347
rect 1678 -397 1744 -381
<< polycont >>
rect -1728 347 -1694 381
rect -1610 347 -1576 381
rect -1492 347 -1458 381
rect -1374 347 -1340 381
rect -1256 347 -1222 381
rect -1138 347 -1104 381
rect -1020 347 -986 381
rect -902 347 -868 381
rect -784 347 -750 381
rect -666 347 -632 381
rect -548 347 -514 381
rect -430 347 -396 381
rect -312 347 -278 381
rect -194 347 -160 381
rect -76 347 -42 381
rect 42 347 76 381
rect 160 347 194 381
rect 278 347 312 381
rect 396 347 430 381
rect 514 347 548 381
rect 632 347 666 381
rect 750 347 784 381
rect 868 347 902 381
rect 986 347 1020 381
rect 1104 347 1138 381
rect 1222 347 1256 381
rect 1340 347 1374 381
rect 1458 347 1492 381
rect 1576 347 1610 381
rect 1694 347 1728 381
rect -1728 -381 -1694 -347
rect -1610 -381 -1576 -347
rect -1492 -381 -1458 -347
rect -1374 -381 -1340 -347
rect -1256 -381 -1222 -347
rect -1138 -381 -1104 -347
rect -1020 -381 -986 -347
rect -902 -381 -868 -347
rect -784 -381 -750 -347
rect -666 -381 -632 -347
rect -548 -381 -514 -347
rect -430 -381 -396 -347
rect -312 -381 -278 -347
rect -194 -381 -160 -347
rect -76 -381 -42 -347
rect 42 -381 76 -347
rect 160 -381 194 -347
rect 278 -381 312 -347
rect 396 -381 430 -347
rect 514 -381 548 -347
rect 632 -381 666 -347
rect 750 -381 784 -347
rect 868 -381 902 -347
rect 986 -381 1020 -347
rect 1104 -381 1138 -347
rect 1222 -381 1256 -347
rect 1340 -381 1374 -347
rect 1458 -381 1492 -347
rect 1576 -381 1610 -347
rect 1694 -381 1728 -347
<< locali >>
rect -1901 449 -1805 483
rect 1805 449 1901 483
rect -1901 387 -1867 449
rect 1867 387 1901 449
rect -1744 347 -1728 381
rect -1694 347 -1678 381
rect -1626 347 -1610 381
rect -1576 347 -1560 381
rect -1508 347 -1492 381
rect -1458 347 -1442 381
rect -1390 347 -1374 381
rect -1340 347 -1324 381
rect -1272 347 -1256 381
rect -1222 347 -1206 381
rect -1154 347 -1138 381
rect -1104 347 -1088 381
rect -1036 347 -1020 381
rect -986 347 -970 381
rect -918 347 -902 381
rect -868 347 -852 381
rect -800 347 -784 381
rect -750 347 -734 381
rect -682 347 -666 381
rect -632 347 -616 381
rect -564 347 -548 381
rect -514 347 -498 381
rect -446 347 -430 381
rect -396 347 -380 381
rect -328 347 -312 381
rect -278 347 -262 381
rect -210 347 -194 381
rect -160 347 -144 381
rect -92 347 -76 381
rect -42 347 -26 381
rect 26 347 42 381
rect 76 347 92 381
rect 144 347 160 381
rect 194 347 210 381
rect 262 347 278 381
rect 312 347 328 381
rect 380 347 396 381
rect 430 347 446 381
rect 498 347 514 381
rect 548 347 564 381
rect 616 347 632 381
rect 666 347 682 381
rect 734 347 750 381
rect 784 347 800 381
rect 852 347 868 381
rect 902 347 918 381
rect 970 347 986 381
rect 1020 347 1036 381
rect 1088 347 1104 381
rect 1138 347 1154 381
rect 1206 347 1222 381
rect 1256 347 1272 381
rect 1324 347 1340 381
rect 1374 347 1390 381
rect 1442 347 1458 381
rect 1492 347 1508 381
rect 1560 347 1576 381
rect 1610 347 1626 381
rect 1678 347 1694 381
rect 1728 347 1744 381
rect -1787 288 -1753 304
rect -1787 -304 -1753 -288
rect -1669 288 -1635 304
rect -1669 -304 -1635 -288
rect -1551 288 -1517 304
rect -1551 -304 -1517 -288
rect -1433 288 -1399 304
rect -1433 -304 -1399 -288
rect -1315 288 -1281 304
rect -1315 -304 -1281 -288
rect -1197 288 -1163 304
rect -1197 -304 -1163 -288
rect -1079 288 -1045 304
rect -1079 -304 -1045 -288
rect -961 288 -927 304
rect -961 -304 -927 -288
rect -843 288 -809 304
rect -843 -304 -809 -288
rect -725 288 -691 304
rect -725 -304 -691 -288
rect -607 288 -573 304
rect -607 -304 -573 -288
rect -489 288 -455 304
rect -489 -304 -455 -288
rect -371 288 -337 304
rect -371 -304 -337 -288
rect -253 288 -219 304
rect -253 -304 -219 -288
rect -135 288 -101 304
rect -135 -304 -101 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 101 288 135 304
rect 101 -304 135 -288
rect 219 288 253 304
rect 219 -304 253 -288
rect 337 288 371 304
rect 337 -304 371 -288
rect 455 288 489 304
rect 455 -304 489 -288
rect 573 288 607 304
rect 573 -304 607 -288
rect 691 288 725 304
rect 691 -304 725 -288
rect 809 288 843 304
rect 809 -304 843 -288
rect 927 288 961 304
rect 927 -304 961 -288
rect 1045 288 1079 304
rect 1045 -304 1079 -288
rect 1163 288 1197 304
rect 1163 -304 1197 -288
rect 1281 288 1315 304
rect 1281 -304 1315 -288
rect 1399 288 1433 304
rect 1399 -304 1433 -288
rect 1517 288 1551 304
rect 1517 -304 1551 -288
rect 1635 288 1669 304
rect 1635 -304 1669 -288
rect 1753 288 1787 304
rect 1753 -304 1787 -288
rect -1744 -381 -1728 -347
rect -1694 -381 -1678 -347
rect -1626 -381 -1610 -347
rect -1576 -381 -1560 -347
rect -1508 -381 -1492 -347
rect -1458 -381 -1442 -347
rect -1390 -381 -1374 -347
rect -1340 -381 -1324 -347
rect -1272 -381 -1256 -347
rect -1222 -381 -1206 -347
rect -1154 -381 -1138 -347
rect -1104 -381 -1088 -347
rect -1036 -381 -1020 -347
rect -986 -381 -970 -347
rect -918 -381 -902 -347
rect -868 -381 -852 -347
rect -800 -381 -784 -347
rect -750 -381 -734 -347
rect -682 -381 -666 -347
rect -632 -381 -616 -347
rect -564 -381 -548 -347
rect -514 -381 -498 -347
rect -446 -381 -430 -347
rect -396 -381 -380 -347
rect -328 -381 -312 -347
rect -278 -381 -262 -347
rect -210 -381 -194 -347
rect -160 -381 -144 -347
rect -92 -381 -76 -347
rect -42 -381 -26 -347
rect 26 -381 42 -347
rect 76 -381 92 -347
rect 144 -381 160 -347
rect 194 -381 210 -347
rect 262 -381 278 -347
rect 312 -381 328 -347
rect 380 -381 396 -347
rect 430 -381 446 -347
rect 498 -381 514 -347
rect 548 -381 564 -347
rect 616 -381 632 -347
rect 666 -381 682 -347
rect 734 -381 750 -347
rect 784 -381 800 -347
rect 852 -381 868 -347
rect 902 -381 918 -347
rect 970 -381 986 -347
rect 1020 -381 1036 -347
rect 1088 -381 1104 -347
rect 1138 -381 1154 -347
rect 1206 -381 1222 -347
rect 1256 -381 1272 -347
rect 1324 -381 1340 -347
rect 1374 -381 1390 -347
rect 1442 -381 1458 -347
rect 1492 -381 1508 -347
rect 1560 -381 1576 -347
rect 1610 -381 1626 -347
rect 1678 -381 1694 -347
rect 1728 -381 1744 -347
rect -1901 -449 -1867 -387
rect 1867 -449 1901 -387
rect -1901 -483 -1805 -449
rect 1805 -483 1901 -449
<< viali >>
rect -1728 347 -1694 381
rect -1610 347 -1576 381
rect -1492 347 -1458 381
rect -1374 347 -1340 381
rect -1256 347 -1222 381
rect -1138 347 -1104 381
rect -1020 347 -986 381
rect -902 347 -868 381
rect -784 347 -750 381
rect -666 347 -632 381
rect -548 347 -514 381
rect -430 347 -396 381
rect -312 347 -278 381
rect -194 347 -160 381
rect -76 347 -42 381
rect 42 347 76 381
rect 160 347 194 381
rect 278 347 312 381
rect 396 347 430 381
rect 514 347 548 381
rect 632 347 666 381
rect 750 347 784 381
rect 868 347 902 381
rect 986 347 1020 381
rect 1104 347 1138 381
rect 1222 347 1256 381
rect 1340 347 1374 381
rect 1458 347 1492 381
rect 1576 347 1610 381
rect 1694 347 1728 381
rect -1787 -288 -1753 288
rect -1669 -288 -1635 288
rect -1551 -288 -1517 288
rect -1433 -288 -1399 288
rect -1315 -288 -1281 288
rect -1197 -288 -1163 288
rect -1079 -288 -1045 288
rect -961 -288 -927 288
rect -843 -288 -809 288
rect -725 -288 -691 288
rect -607 -288 -573 288
rect -489 -288 -455 288
rect -371 -288 -337 288
rect -253 -288 -219 288
rect -135 -288 -101 288
rect -17 -288 17 288
rect 101 -288 135 288
rect 219 -288 253 288
rect 337 -288 371 288
rect 455 -288 489 288
rect 573 -288 607 288
rect 691 -288 725 288
rect 809 -288 843 288
rect 927 -288 961 288
rect 1045 -288 1079 288
rect 1163 -288 1197 288
rect 1281 -288 1315 288
rect 1399 -288 1433 288
rect 1517 -288 1551 288
rect 1635 -288 1669 288
rect 1753 -288 1787 288
rect -1728 -381 -1694 -347
rect -1610 -381 -1576 -347
rect -1492 -381 -1458 -347
rect -1374 -381 -1340 -347
rect -1256 -381 -1222 -347
rect -1138 -381 -1104 -347
rect -1020 -381 -986 -347
rect -902 -381 -868 -347
rect -784 -381 -750 -347
rect -666 -381 -632 -347
rect -548 -381 -514 -347
rect -430 -381 -396 -347
rect -312 -381 -278 -347
rect -194 -381 -160 -347
rect -76 -381 -42 -347
rect 42 -381 76 -347
rect 160 -381 194 -347
rect 278 -381 312 -347
rect 396 -381 430 -347
rect 514 -381 548 -347
rect 632 -381 666 -347
rect 750 -381 784 -347
rect 868 -381 902 -347
rect 986 -381 1020 -347
rect 1104 -381 1138 -347
rect 1222 -381 1256 -347
rect 1340 -381 1374 -347
rect 1458 -381 1492 -347
rect 1576 -381 1610 -347
rect 1694 -381 1728 -347
<< metal1 >>
rect -1740 381 -1682 387
rect -1740 347 -1728 381
rect -1694 347 -1682 381
rect -1740 341 -1682 347
rect -1622 381 -1564 387
rect -1622 347 -1610 381
rect -1576 347 -1564 381
rect -1622 341 -1564 347
rect -1504 381 -1446 387
rect -1504 347 -1492 381
rect -1458 347 -1446 381
rect -1504 341 -1446 347
rect -1386 381 -1328 387
rect -1386 347 -1374 381
rect -1340 347 -1328 381
rect -1386 341 -1328 347
rect -1268 381 -1210 387
rect -1268 347 -1256 381
rect -1222 347 -1210 381
rect -1268 341 -1210 347
rect -1150 381 -1092 387
rect -1150 347 -1138 381
rect -1104 347 -1092 381
rect -1150 341 -1092 347
rect -1032 381 -974 387
rect -1032 347 -1020 381
rect -986 347 -974 381
rect -1032 341 -974 347
rect -914 381 -856 387
rect -914 347 -902 381
rect -868 347 -856 381
rect -914 341 -856 347
rect -796 381 -738 387
rect -796 347 -784 381
rect -750 347 -738 381
rect -796 341 -738 347
rect -678 381 -620 387
rect -678 347 -666 381
rect -632 347 -620 381
rect -678 341 -620 347
rect -560 381 -502 387
rect -560 347 -548 381
rect -514 347 -502 381
rect -560 341 -502 347
rect -442 381 -384 387
rect -442 347 -430 381
rect -396 347 -384 381
rect -442 341 -384 347
rect -324 381 -266 387
rect -324 347 -312 381
rect -278 347 -266 381
rect -324 341 -266 347
rect -206 381 -148 387
rect -206 347 -194 381
rect -160 347 -148 381
rect -206 341 -148 347
rect -88 381 -30 387
rect -88 347 -76 381
rect -42 347 -30 381
rect -88 341 -30 347
rect 30 381 88 387
rect 30 347 42 381
rect 76 347 88 381
rect 30 341 88 347
rect 148 381 206 387
rect 148 347 160 381
rect 194 347 206 381
rect 148 341 206 347
rect 266 381 324 387
rect 266 347 278 381
rect 312 347 324 381
rect 266 341 324 347
rect 384 381 442 387
rect 384 347 396 381
rect 430 347 442 381
rect 384 341 442 347
rect 502 381 560 387
rect 502 347 514 381
rect 548 347 560 381
rect 502 341 560 347
rect 620 381 678 387
rect 620 347 632 381
rect 666 347 678 381
rect 620 341 678 347
rect 738 381 796 387
rect 738 347 750 381
rect 784 347 796 381
rect 738 341 796 347
rect 856 381 914 387
rect 856 347 868 381
rect 902 347 914 381
rect 856 341 914 347
rect 974 381 1032 387
rect 974 347 986 381
rect 1020 347 1032 381
rect 974 341 1032 347
rect 1092 381 1150 387
rect 1092 347 1104 381
rect 1138 347 1150 381
rect 1092 341 1150 347
rect 1210 381 1268 387
rect 1210 347 1222 381
rect 1256 347 1268 381
rect 1210 341 1268 347
rect 1328 381 1386 387
rect 1328 347 1340 381
rect 1374 347 1386 381
rect 1328 341 1386 347
rect 1446 381 1504 387
rect 1446 347 1458 381
rect 1492 347 1504 381
rect 1446 341 1504 347
rect 1564 381 1622 387
rect 1564 347 1576 381
rect 1610 347 1622 381
rect 1564 341 1622 347
rect 1682 381 1740 387
rect 1682 347 1694 381
rect 1728 347 1740 381
rect 1682 341 1740 347
rect -1793 288 -1747 300
rect -1793 -288 -1787 288
rect -1753 -288 -1747 288
rect -1793 -300 -1747 -288
rect -1675 288 -1629 300
rect -1675 -288 -1669 288
rect -1635 -288 -1629 288
rect -1675 -300 -1629 -288
rect -1557 288 -1511 300
rect -1557 -288 -1551 288
rect -1517 -288 -1511 288
rect -1557 -300 -1511 -288
rect -1439 288 -1393 300
rect -1439 -288 -1433 288
rect -1399 -288 -1393 288
rect -1439 -300 -1393 -288
rect -1321 288 -1275 300
rect -1321 -288 -1315 288
rect -1281 -288 -1275 288
rect -1321 -300 -1275 -288
rect -1203 288 -1157 300
rect -1203 -288 -1197 288
rect -1163 -288 -1157 288
rect -1203 -300 -1157 -288
rect -1085 288 -1039 300
rect -1085 -288 -1079 288
rect -1045 -288 -1039 288
rect -1085 -300 -1039 -288
rect -967 288 -921 300
rect -967 -288 -961 288
rect -927 -288 -921 288
rect -967 -300 -921 -288
rect -849 288 -803 300
rect -849 -288 -843 288
rect -809 -288 -803 288
rect -849 -300 -803 -288
rect -731 288 -685 300
rect -731 -288 -725 288
rect -691 -288 -685 288
rect -731 -300 -685 -288
rect -613 288 -567 300
rect -613 -288 -607 288
rect -573 -288 -567 288
rect -613 -300 -567 -288
rect -495 288 -449 300
rect -495 -288 -489 288
rect -455 -288 -449 288
rect -495 -300 -449 -288
rect -377 288 -331 300
rect -377 -288 -371 288
rect -337 -288 -331 288
rect -377 -300 -331 -288
rect -259 288 -213 300
rect -259 -288 -253 288
rect -219 -288 -213 288
rect -259 -300 -213 -288
rect -141 288 -95 300
rect -141 -288 -135 288
rect -101 -288 -95 288
rect -141 -300 -95 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 95 288 141 300
rect 95 -288 101 288
rect 135 -288 141 288
rect 95 -300 141 -288
rect 213 288 259 300
rect 213 -288 219 288
rect 253 -288 259 288
rect 213 -300 259 -288
rect 331 288 377 300
rect 331 -288 337 288
rect 371 -288 377 288
rect 331 -300 377 -288
rect 449 288 495 300
rect 449 -288 455 288
rect 489 -288 495 288
rect 449 -300 495 -288
rect 567 288 613 300
rect 567 -288 573 288
rect 607 -288 613 288
rect 567 -300 613 -288
rect 685 288 731 300
rect 685 -288 691 288
rect 725 -288 731 288
rect 685 -300 731 -288
rect 803 288 849 300
rect 803 -288 809 288
rect 843 -288 849 288
rect 803 -300 849 -288
rect 921 288 967 300
rect 921 -288 927 288
rect 961 -288 967 288
rect 921 -300 967 -288
rect 1039 288 1085 300
rect 1039 -288 1045 288
rect 1079 -288 1085 288
rect 1039 -300 1085 -288
rect 1157 288 1203 300
rect 1157 -288 1163 288
rect 1197 -288 1203 288
rect 1157 -300 1203 -288
rect 1275 288 1321 300
rect 1275 -288 1281 288
rect 1315 -288 1321 288
rect 1275 -300 1321 -288
rect 1393 288 1439 300
rect 1393 -288 1399 288
rect 1433 -288 1439 288
rect 1393 -300 1439 -288
rect 1511 288 1557 300
rect 1511 -288 1517 288
rect 1551 -288 1557 288
rect 1511 -300 1557 -288
rect 1629 288 1675 300
rect 1629 -288 1635 288
rect 1669 -288 1675 288
rect 1629 -300 1675 -288
rect 1747 288 1793 300
rect 1747 -288 1753 288
rect 1787 -288 1793 288
rect 1747 -300 1793 -288
rect -1740 -347 -1682 -341
rect -1740 -381 -1728 -347
rect -1694 -381 -1682 -347
rect -1740 -387 -1682 -381
rect -1622 -347 -1564 -341
rect -1622 -381 -1610 -347
rect -1576 -381 -1564 -347
rect -1622 -387 -1564 -381
rect -1504 -347 -1446 -341
rect -1504 -381 -1492 -347
rect -1458 -381 -1446 -347
rect -1504 -387 -1446 -381
rect -1386 -347 -1328 -341
rect -1386 -381 -1374 -347
rect -1340 -381 -1328 -347
rect -1386 -387 -1328 -381
rect -1268 -347 -1210 -341
rect -1268 -381 -1256 -347
rect -1222 -381 -1210 -347
rect -1268 -387 -1210 -381
rect -1150 -347 -1092 -341
rect -1150 -381 -1138 -347
rect -1104 -381 -1092 -347
rect -1150 -387 -1092 -381
rect -1032 -347 -974 -341
rect -1032 -381 -1020 -347
rect -986 -381 -974 -347
rect -1032 -387 -974 -381
rect -914 -347 -856 -341
rect -914 -381 -902 -347
rect -868 -381 -856 -347
rect -914 -387 -856 -381
rect -796 -347 -738 -341
rect -796 -381 -784 -347
rect -750 -381 -738 -347
rect -796 -387 -738 -381
rect -678 -347 -620 -341
rect -678 -381 -666 -347
rect -632 -381 -620 -347
rect -678 -387 -620 -381
rect -560 -347 -502 -341
rect -560 -381 -548 -347
rect -514 -381 -502 -347
rect -560 -387 -502 -381
rect -442 -347 -384 -341
rect -442 -381 -430 -347
rect -396 -381 -384 -347
rect -442 -387 -384 -381
rect -324 -347 -266 -341
rect -324 -381 -312 -347
rect -278 -381 -266 -347
rect -324 -387 -266 -381
rect -206 -347 -148 -341
rect -206 -381 -194 -347
rect -160 -381 -148 -347
rect -206 -387 -148 -381
rect -88 -347 -30 -341
rect -88 -381 -76 -347
rect -42 -381 -30 -347
rect -88 -387 -30 -381
rect 30 -347 88 -341
rect 30 -381 42 -347
rect 76 -381 88 -347
rect 30 -387 88 -381
rect 148 -347 206 -341
rect 148 -381 160 -347
rect 194 -381 206 -347
rect 148 -387 206 -381
rect 266 -347 324 -341
rect 266 -381 278 -347
rect 312 -381 324 -347
rect 266 -387 324 -381
rect 384 -347 442 -341
rect 384 -381 396 -347
rect 430 -381 442 -347
rect 384 -387 442 -381
rect 502 -347 560 -341
rect 502 -381 514 -347
rect 548 -381 560 -347
rect 502 -387 560 -381
rect 620 -347 678 -341
rect 620 -381 632 -347
rect 666 -381 678 -347
rect 620 -387 678 -381
rect 738 -347 796 -341
rect 738 -381 750 -347
rect 784 -381 796 -347
rect 738 -387 796 -381
rect 856 -347 914 -341
rect 856 -381 868 -347
rect 902 -381 914 -347
rect 856 -387 914 -381
rect 974 -347 1032 -341
rect 974 -381 986 -347
rect 1020 -381 1032 -347
rect 974 -387 1032 -381
rect 1092 -347 1150 -341
rect 1092 -381 1104 -347
rect 1138 -381 1150 -347
rect 1092 -387 1150 -381
rect 1210 -347 1268 -341
rect 1210 -381 1222 -347
rect 1256 -381 1268 -347
rect 1210 -387 1268 -381
rect 1328 -347 1386 -341
rect 1328 -381 1340 -347
rect 1374 -381 1386 -347
rect 1328 -387 1386 -381
rect 1446 -347 1504 -341
rect 1446 -381 1458 -347
rect 1492 -381 1504 -347
rect 1446 -387 1504 -381
rect 1564 -347 1622 -341
rect 1564 -381 1576 -347
rect 1610 -381 1622 -347
rect 1564 -387 1622 -381
rect 1682 -347 1740 -341
rect 1682 -381 1694 -347
rect 1728 -381 1740 -347
rect 1682 -387 1740 -381
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1884 -466 1884 466
string parameters w 3 l 0.3 m 1 nf 30 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
